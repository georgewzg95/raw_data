//////////////////////////////////////////////////////////////////////////////////
// Company:         
// Engineer:        IK
// 
// Design Name:
// Module Name:
// Project Name:    PowerOnReset Module
// Target Devices:  

// Description: 
//
//
// Revision: 
// Revision 0.01 - File Created
//
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module por_module #(parameter p_LEN = 0)
(
    // SYS_CON
    input           i_clk,
    // POR out
    output  reg     o_por
);
//////////////////////////////////////////////////////////////////////////////////
    // por-cnt
    reg [p_LEN-1:0]   sv_por_cnt=0;
    
//////////////////////////////////////////////////////////////////////////////////
//
// PowerOnReset logic
//
always @ (posedge i_clk)
begin   :   POR_LOGIC
    // inner
    if (!sv_por_cnt[p_LEN-1])
        sv_por_cnt <= sv_por_cnt + 1'b1;
    // out
    o_por <= !sv_por_cnt[p_LEN-1];
end
//////////////////////////////////////////////////////////////////////////////////
endmodule

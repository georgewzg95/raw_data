//////////////////////////////////////////////////////////////////////////////////
// Company:         
// Engineer:        IK
// 
// Create Date:     
// Design Name:     
// Module Name:     clk_module
// Project Name:    
// Target Devices:  
// Tool versions:   
// Description:     
//                  
//                  
// Revision: 
// Revision 0.01 - File Created, 
//
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module rst_sync
(
    // SYS_CON
    input       i_clk,
    // iRST
    input       i_arst,
    // oRST
    output      o_srst
);
//////////////////////////////////////////////////////////////////////////////////
// ??
localparam  lp_RW = 4;
//////////////////////////////////////////////////////////////////////////////////
    // sync-rst-chain
    reg     [lp_RW-1:0]   sv_srst;
//////////////////////////////////////////////////////////////////////////////////
    // oRST
    assign o_srst = !sv_srst[lp_RW-1];
//////////////////////////////////////////////////////////////////////////////////
//
// ??
//
always @ (posedge i_clk or posedge i_arst)
begin   :   SRST_LOGIC
    if (i_arst)
        sv_srst <= 0;
    else
        sv_srst <= {sv_srst[2:0], 1'b1};
end
//////////////////////////////////////////////////////////////////////////////////
endmodule

//-------------------------------------------------------------------------
//
// File name    :  ldpc_cn.v
// Title        :
//              :
// Purpose      : Check node holder/message calculator.  Stores the sign
//              : of each received message, along with
//
// ----------------------------------------------------------------------
// Revision History :
// ----------------------------------------------------------------------
//   Ver  :| Author   :| Mod. Date   :| Changes Made:
//   v1.0  | JTC      :| 2008/07/02  :|
// ----------------------------------------------------------------------
`timescale 1ns/10ps

module ldpc_cn #(
  parameter FOLDFACTOR     = 1,
  parameter LLRWIDTH       = 6
)(
  input clk,
  input rst,

  // clear RAM iteration count at start-up
  input      llr_access,
  input[7:0] llr_addr,
  input      llr_din_we,

  // message I/O
  input                   iteration,         // toggle each iteration
  input                   first_half,
  input                   first_iteration,   // don't need to subtract-off previous message!
  input                   cn_we,
  input                   cn_rd,
  input                   disable_cn, // parity mix disables one node
  input[7+FOLDFACTOR-1:0] addr_cn,
  input[LLRWIDTH-1:0]     sh_msg,
  output[LLRWIDTH-1:0]    cn_msg,

  // Attached MSG RAM, 135xMSG_WIDTH
  output                         dnmsg_we,
  output[7+FOLDFACTOR-1:0]       dnmsg_wraddr,
  output[7+FOLDFACTOR-1:0]       dnmsg_rdaddr,
  output[17+4*(LLRWIDTH-1)+31:0] dnmsg_din,
  input[17+4*(LLRWIDTH-1)+31:0]  dnmsg_dout
);

// Detect illegal writes
// synthesis translate_off
integer accesses[0:5];
reg     a_run;
integer temp_loopvar;

always @( posedge rst, posedge clk )
  if( rst )
    for( temp_loopvar=0; temp_loopvar<6; temp_loopvar=temp_loopvar+1 )
      accesses[temp_loopvar] = -1;
  else
  begin
    for( temp_loopvar=5; temp_loopvar>0; temp_loopvar=temp_loopvar-1 )
    begin
      accesses[temp_loopvar] = accesses[temp_loopvar-1];
      if( !(cn_we|cn_rd) )
        accesses[0] = -1;
      else
        accesses[0] = addr_cn;
    end
    
    a_run = 1;
    
    for( temp_loopvar=1; temp_loopvar<6; temp_loopvar=temp_loopvar+1 )
    begin
      a_run = a_run & (accesses[temp_loopvar]==addr_cn);
      if( !a_run && (cn_we|cn_rd) && (accesses[temp_loopvar]==addr_cn) )
        $display( "%0t: Bad access, addresses %0d", $time(), addr_cn );
     end
  end
// synthesis translate_on

assign dnmsg_rdaddr = llr_access ? llr_addr : addr_cn;

/***********************************
 * Calc message/update message RAM *
 * Combine 1's complement numbers  *
 * Saturate to one bit fewer than  *
 * input width                     *
 ***********************************/
function[LLRWIDTH-1:0] SubSaturate( input[LLRWIDTH-1:0] a,
                                    input[LLRWIDTH-1:0] b );
  reg[LLRWIDTH-1:0] sum;
  reg[LLRWIDTH-2:0] diffa;
  reg[LLRWIDTH-2:0] diffb;
  reg[LLRWIDTH-3:0] sat_sum;
  reg[LLRWIDTH-3:0] sat_diffa;
  reg[LLRWIDTH-3:0] sat_diffb;
  reg               add;
  reg               b_big;
  reg               sign;
  reg[LLRWIDTH-1:0] result;
begin
  // basic calculations
  sum   = {1'b0, a[LLRWIDTH-2:0]} + {1'b0, b[LLRWIDTH-2:0]};
  diffa = a[LLRWIDTH-2:0] - b[LLRWIDTH-2:0];
  diffb = b[LLRWIDTH-2:0] - a[LLRWIDTH-2:0];

  // saturate
  if( sum[LLRWIDTH-1:LLRWIDTH-2]!=2'b00  )
    sat_sum = { (LLRWIDTH-2){1'b1} };
  else
    sat_sum = sum[LLRWIDTH-3:0];

  if( diffa[LLRWIDTH-2]  )
    sat_diffa = { (LLRWIDTH-2){1'b1} };
  else
    sat_diffa = diffa[LLRWIDTH-3:0];

  if( diffb[LLRWIDTH-2]  )
    sat_diffb = { (LLRWIDTH-2){1'b1} };
  else
    sat_diffb = diffb[LLRWIDTH-3:0];

  // control bits
  add   = a[LLRWIDTH-1]!=b[LLRWIDTH-1];
  b_big = a[LLRWIDTH-2:0]<b[LLRWIDTH-2:0];
  sign  = b_big ? ~b[LLRWIDTH-1] : a[LLRWIDTH-1];

  if( add )
    result = { sign, 1'b0, sat_sum };
  else if( b_big )
    result = { sign, 1'b0, sat_diffb };
  else
    result = { sign, 1'b0, sat_diffa };

  SubSaturate = result;
end
endfunction

/**************************************
 * Align some signals with RAM output *
 **************************************/
localparam RAM_LATENCY = 2;

integer loopvar1;

reg                   cn_rd_del[0:RAM_LATENCY-1];
reg                   cn_we_del[0:RAM_LATENCY-1];
reg[LLRWIDTH-1:0]     sh_msg_del[0:RAM_LATENCY-1];
reg[7+FOLDFACTOR-1:0] addr_cn_del[0:RAM_LATENCY-1];

reg repeat_access;

wire                   cn_rd_aligned_ram;
wire                   cn_we_aligned_ram;
wire[LLRWIDTH-1:0]     sh_msg_aligned_ram;
wire[7+FOLDFACTOR-1:0] addr_cn_aligned_ram;

assign cn_rd_aligned_ram   = cn_rd_del[RAM_LATENCY-1];
assign cn_we_aligned_ram   = cn_we_del[RAM_LATENCY-1];
assign sh_msg_aligned_ram  = sh_msg_del[RAM_LATENCY-1];
assign addr_cn_aligned_ram = addr_cn_del[RAM_LATENCY-1];

always @( posedge rst, posedge clk )
  if( rst )
  begin
    for( loopvar1=0; loopvar1<RAM_LATENCY; loopvar1=loopvar1+1 )
    begin
      cn_rd_del[loopvar1]   <= 0;
      cn_we_del[loopvar1]   <= 0;
      sh_msg_del[loopvar1]  <= 0;
      addr_cn_del[loopvar1] <= 0;
    end
    repeat_access <= 0;
  end
  else
  begin
    cn_rd_del[0]   <= cn_rd & ~disable_cn;
    cn_we_del[0]   <= cn_we & ~disable_cn;
    sh_msg_del[0]  <= sh_msg;
    addr_cn_del[0] <= addr_cn;

    for( loopvar1=1; loopvar1<RAM_LATENCY; loopvar1=loopvar1+1 )
    begin
      cn_rd_del[loopvar1]   <= cn_rd_del[loopvar1 -1];
      cn_we_del[loopvar1]   <= cn_we_del[loopvar1 -1];
      sh_msg_del[loopvar1]  <= sh_msg_del[loopvar1 -1];
      addr_cn_del[loopvar1] <= addr_cn_del[loopvar1 -1];
    end

    repeat_access <= (addr_cn_del[RAM_LATENCY-1]==addr_cn_del[RAM_LATENCY-2]) &&
                     ((cn_we_del[RAM_LATENCY-1] && cn_we_del[RAM_LATENCY-2]) ||
                      (cn_rd_del[RAM_LATENCY-1] && cn_rd_del[RAM_LATENCY-2]));
  end

/****************************
 * Pipe stage 0:            *
 * Register bits out of RAM *
 ****************************/
wire start_over;
wire switch_up;

reg[4:0]          old_leastpos;
reg[4:0]          old_last_leastpos;
reg               old_sign_result;
reg[4:0]          old_count;
reg[LLRWIDTH-2:0] old_least_llr;
reg[LLRWIDTH-2:0] old_nextleast_llr;
reg[LLRWIDTH-2:0] old_last_least_llr;
reg[LLRWIDTH-2:0] old_last_nextleast_llr;
reg               old_last_sign_result;
reg[29:0]         old_signs;

reg[LLRWIDTH-1:0] sh_msg_aligned_old;
reg               start_over_aligned_old;
reg               repeat_access_aligned_old;
reg               cn_we_aligned_old;

// restart calculations and count if RAM's iteration != controller's iteration
assign start_over = (iteration!=dnmsg_dout[0]) & !repeat_access;

// restart count when switching from downstream to upstream messages
assign switch_up  = ~first_half & ~dnmsg_dout[1] & !repeat_access;

always @( posedge clk, posedge rst )
  if( rst )
  begin
    old_count                 <= 0;
    old_leastpos              <= 0;
    old_last_leastpos         <= 0;
    old_sign_result           <= 0;
    old_least_llr             <= 0;
    old_nextleast_llr         <= 0;
    old_last_least_llr        <= 0;
    old_last_nextleast_llr    <= 0;
    old_last_sign_result      <= 0;
    old_signs                 <= 0;
    sh_msg_aligned_old        <= 0;
    start_over_aligned_old    <= 0;
    cn_we_aligned_old         <= 0;
    repeat_access_aligned_old <= 0;
  end
  else
  begin
    if( repeat_access )
      old_count <= old_count + 1;
    else
      old_count <= (start_over | switch_up) ? 0 : dnmsg_dout[16:12];

    old_leastpos           <= dnmsg_dout[6:2];
    old_last_leastpos      <= dnmsg_dout[11:7];
    old_least_llr          <= dnmsg_dout[16 +1*(LLRWIDTH-1) -: LLRWIDTH-1];
    old_nextleast_llr      <= dnmsg_dout[16 +2*(LLRWIDTH-1) -: LLRWIDTH-1];
    old_last_least_llr     <= dnmsg_dout[16 +3*(LLRWIDTH-1) -: LLRWIDTH-1];
    old_last_nextleast_llr <= dnmsg_dout[16 +4*(LLRWIDTH-1) -: LLRWIDTH-1];
    old_sign_result        <= dnmsg_dout[16 +4*(LLRWIDTH-1)+1];
    old_last_sign_result   <= dnmsg_dout[16 +4*(LLRWIDTH-1)+2];
    old_signs              <= dnmsg_dout[16 +4*(LLRWIDTH-1)+32 -: 30];

    sh_msg_aligned_old        <= sh_msg_aligned_ram;
    start_over_aligned_old    <= start_over;
    cn_we_aligned_old         <= cn_we_aligned_ram;
    repeat_access_aligned_old <= repeat_access;
  end

/***************************
 * Pipe 1a:                *
 * Create outgoing message *
 ***************************/
reg[LLRWIDTH-1:0] cn_msg_int;

assign cn_msg = cn_msg_int;

always @( posedge rst, posedge clk )
  if( rst )
    cn_msg_int <= 0;
  else
  begin
    // sign val
    cn_msg_int[LLRWIDTH-1] <= old_sign_result ^ old_signs[old_count];

    // min result
    if( old_count==old_leastpos )
      cn_msg_int[LLRWIDTH-2:0] <= old_nextleast_llr;
    else
      cn_msg_int[LLRWIDTH-2:0] <= old_least_llr;
  end

/****************************************************************
 * Pipe stage 1b:                                               *
 * Calculate fixed_msg = downlink message - last uplink message *
 ****************************************************************/
wire[LLRWIDTH-1:0] offset_val;
reg[LLRWIDTH-1:0]  fixed_msg;

reg[LLRWIDTH-2:0] old_least_llr_del;
reg[LLRWIDTH-2:0] old_nextleast_llr_del;
reg[4:0]          old_count_del;
reg[4:0]          old_leastpos_del;
reg[29:0]         old_signs_del;
reg               old_sign_result_del;
reg               old_last_sign_result_del;
reg[4:0]          old_last_leastpos_del;
reg[LLRWIDTH-2:0] old_last_least_llr_del;
reg[LLRWIDTH-2:0] old_last_nextleast_llr_del;

reg start_over_aligned_msg;
reg cn_we_aligned_msg;
reg repeat_access_aligned_msg;

assign offset_val = first_iteration ? 0
                      : (old_count==old_last_leastpos) ? { old_last_sign_result^old_signs[old_count], old_last_nextleast_llr }
                        : { old_last_sign_result^old_signs[old_count], old_last_least_llr };

always @( posedge rst, posedge clk )
  if( rst )
  begin
    fixed_msg                  <= 0;
    old_least_llr_del          <= 0;
    old_nextleast_llr_del      <= 0;
    old_count_del              <= 0;
    old_leastpos_del           <= 0;
    old_signs_del              <= 0;
    old_sign_result_del        <= 0;
    old_last_sign_result_del   <= 0;
    old_last_leastpos_del      <= 0;
    old_last_least_llr_del     <= 0;
    old_last_nextleast_llr_del <= 0;
    start_over_aligned_msg     <= 0;
    cn_we_aligned_msg          <= 0;
    repeat_access_aligned_msg  <= 0;
  end
  else
  begin
    fixed_msg <= SubSaturate( sh_msg_aligned_old, offset_val );

    old_least_llr_del     <= old_least_llr;
    old_nextleast_llr_del <= old_nextleast_llr;
    old_leastpos_del      <= old_leastpos;
    old_signs_del         <= old_signs;
    old_sign_result_del   <= old_sign_result;
    
    old_last_sign_result_del   <= old_last_sign_result;
    old_last_leastpos_del      <= old_last_leastpos;
    old_last_least_llr_del     <= old_last_least_llr;
    old_last_nextleast_llr_del <= old_last_nextleast_llr;

    old_count_del <= old_count;

    start_over_aligned_msg    <= start_over_aligned_old;
    cn_we_aligned_msg         <= cn_we_aligned_old;
    repeat_access_aligned_msg <= repeat_access_aligned_old;
  end

/*******************************************
 * Pipe stage 2:                           *
 * Calculate new values for RAM write-back *
 *******************************************/
reg               new_iteration;
reg               new_up;
reg[4:0]          new_leastpos;
reg               new_last_sign_result;
reg[4:0]          new_last_leastpos;
reg[29:0]         new_signs;
reg               new_sign_result;
reg[4:0]          new_count;
reg[LLRWIDTH-2:0] new_least_llr;
reg[LLRWIDTH-2:0] new_nextleast_llr;
reg[LLRWIDTH-2:0] new_last_least_llr;
reg[LLRWIDTH-2:0] new_last_nextleast_llr;

wire[LLRWIDTH-2:0] muxed_least_llr;
wire[LLRWIDTH-2:0] muxed_nextleast_llr;
wire new_winner;
wire new_2nd;

assign muxed_least_llr     = repeat_access_aligned_msg ? new_least_llr[LLRWIDTH-2:0]
                                                       : old_least_llr_del[LLRWIDTH-2:0];
assign muxed_nextleast_llr = repeat_access_aligned_msg ? new_nextleast_llr[LLRWIDTH-2:0]
                                                       : old_nextleast_llr_del[LLRWIDTH-2:0];

assign new_winner = (fixed_msg[LLRWIDTH-2:0] < muxed_least_llr[LLRWIDTH-2:0]);
assign new_2nd    = ((fixed_msg[LLRWIDTH-2:0] <= muxed_nextleast_llr[LLRWIDTH-2:0])
                      & ~new_winner);

always @( posedge rst, posedge clk )
  if( rst )
  begin
    new_iteration          <= 0;
    new_up                 <= 0;
    new_count              <= 0;
    new_leastpos           <= 0;
    new_least_llr          <= 0;
    new_nextleast_llr      <= 0;
    new_signs              <= 0;
    new_sign_result        <= 0;
    new_last_sign_result   <= 0;
    new_last_leastpos      <= 0;
    new_last_least_llr     <= 0;
    new_last_nextleast_llr <= 0;
  end
  else
  begin
    new_iteration <= iteration | llr_din_we;
    new_up        <= ~first_half;
    new_count     <= old_count_del + 1;

    // assign new smallest LLR
    if( !repeat_access_aligned_msg )
    begin
      new_signs         <= old_signs_del;
      new_leastpos      <= old_leastpos_del;
      new_least_llr     <= old_least_llr_del;
      new_nextleast_llr <= old_nextleast_llr_del;
      new_sign_result   <= old_sign_result_del;
    end

    if( cn_we_aligned_msg )
    begin
      // note: only assigning one bit - others stay at old value
      new_signs[old_count_del] <= fixed_msg[LLRWIDTH-1];

      if( new_winner | start_over_aligned_msg )
      begin
        new_leastpos  <= old_count_del;
        new_least_llr <= fixed_msg[LLRWIDTH-2:0];
      end

      if( start_over_aligned_msg )
        new_nextleast_llr <= { (LLRWIDTH-1){1'b1} };
      else if( new_winner && repeat_access_aligned_msg )
        new_nextleast_llr <= new_least_llr;
      else if( new_winner )
        new_nextleast_llr <= old_least_llr_del;
      else if( new_2nd )
        new_nextleast_llr <= fixed_msg[LLRWIDTH-2:0];

      if( start_over_aligned_msg )
        new_sign_result <= fixed_msg[LLRWIDTH-1];
      else if( repeat_access_aligned_msg )
        new_sign_result <= new_sign_result ^ fixed_msg[LLRWIDTH-1];
      else
        new_sign_result <= old_sign_result_del ^ fixed_msg[LLRWIDTH-1];
    end

    // store old downstream results during upstream messages
    new_last_sign_result   <= first_half ? old_last_sign_result_del   : old_sign_result_del;
    new_last_leastpos      <= first_half ? old_last_leastpos_del      : old_leastpos_del;
    new_last_least_llr     <= first_half ? old_last_least_llr_del     : old_least_llr_del;
    new_last_nextleast_llr <= first_half ? old_last_nextleast_llr_del : old_nextleast_llr_del;
  end

assign dnmsg_din[0]                                = new_iteration;
assign dnmsg_din[1]                                = new_up;
assign dnmsg_din[6:2]                              = new_leastpos;
assign dnmsg_din[11:7]                             = new_last_leastpos;
assign dnmsg_din[16:12]                            = new_count;
assign dnmsg_din[16+ 1*(LLRWIDTH-1) -: LLRWIDTH-1] = new_least_llr;
assign dnmsg_din[16+ 2*(LLRWIDTH-1) -: LLRWIDTH-1] = new_nextleast_llr;
assign dnmsg_din[16+ 3*(LLRWIDTH-1) -: LLRWIDTH-1] = new_last_least_llr;
assign dnmsg_din[16+ 4*(LLRWIDTH-1) -: LLRWIDTH-1] = new_last_nextleast_llr;
assign dnmsg_din[16+ 4*(LLRWIDTH-1) +1]            = new_sign_result;
assign dnmsg_din[16+ 4*(LLRWIDTH-1) +2]            = new_last_sign_result;
assign dnmsg_din[16+ 4*(LLRWIDTH-1) +32 -: 30]     = new_signs;

/******************************************
 * Align some signals with new RAM inputs *
 ******************************************/
localparam CALC_LATENCY = 3;

integer loopvar2;

reg                   we_del2[0:CALC_LATENCY-1];
reg[7+FOLDFACTOR-1:0] addr_del2[0:CALC_LATENCY-1];

assign dnmsg_we     = ~we_del2[CALC_LATENCY -1];
assign dnmsg_wraddr = addr_del2[CALC_LATENCY -1];

always @( posedge clk, posedge rst )
  if( rst )
    for( loopvar2=0; loopvar2<CALC_LATENCY; loopvar2=loopvar2+1 )
    begin
      we_del2[loopvar2]   <= 0;
      addr_del2[loopvar2] <= 0;
    end
  else
  begin
    we_del2[0]   <= cn_we_aligned_ram | cn_rd_aligned_ram;
    addr_del2[0] <= addr_cn_aligned_ram;

    for( loopvar2=1; loopvar2<CALC_LATENCY; loopvar2=loopvar2+1 )
    begin
      we_del2[loopvar2]   <= we_del2[loopvar2 -1];
      addr_del2[loopvar2] <= addr_del2[loopvar2 -1];
    end

    // last stage - mux in LLR values (if CALC_LATENCY=2, this stage
    // supercedes the entire for-loop, above)
    we_del2[CALC_LATENCY-1] <= llr_din_we | we_del2[CALC_LATENCY-2];

    if( llr_din_we )
      addr_del2[CALC_LATENCY-1] <= llr_addr;
    else
      addr_del2[CALC_LATENCY-1] <= addr_del2[CALC_LATENCY-2];
  end

endmodule
//-------------------------------------------------------------------------
//
// File name    :  ldpc_edgetable.v
// Title        :
//              :
// Purpose      : ROM, holds DVB-S2 edge table
//              : Format:
//              : Code pointer: points to the beginning of a code group
//              :   address[12:0]
//              :
//              : Line descriptor : describes the group of parity
//              :                   descriptors that follow
//              :   bits 13:9: # of parity descriptors in this group
//              :   bit 8: indicate that this is the last group of
//              :          parity descriptors for this code group
//              :   bits 7:0: q value for this group
//              : 
//              : Parity descriptor
//              :   bits 15:9: parity location/q, indicates the distance
//              :              to shift VN input to align with CN
//              :   bits 8:0: parity location MOD q, indicates the CN
//              :             address for this check node
//
// ----------------------------------------------------------------------
// Revision History :
// ----------------------------------------------------------------------
//   Ver  :| Author   :| Mod. Date   :| Changes Made:
//   v1.0  | JTC      :| 2008/07/02  :|
// ----------------------------------------------------------------------
`timescale 1ns/10ps

module ldpc_edgetable(
  input        clk,
  input        rst,
  input[12:0]  romaddr,
  output[16:0] romdata
);

reg[16:0] romdata_int;

assign romdata = romdata_int;

always @( posedge rst, posedge clk )
  if( rst )
    romdata_int <= 0;
  else
  case( romaddr )
    0: romdata_int  <= 'h15;   // Code pointer for 1_4
    1: romdata_int  <= 'h150;  // Code pointer for 1_3
    2: romdata_int  <= 'h2f4;  // Code pointer for 2_5
    3: romdata_int  <= 'h4ec;  // Code pointer for 1_2
    4: romdata_int  <= 'h708;  // Code pointer for 3_5
    5: romdata_int  <= 'h9fc;  // Code pointer for 2_3
    6: romdata_int  <= 'hc54;  // Code pointer for 3_4
    7: romdata_int  <= 'hef7;  // Code pointer for 4_5
    8: romdata_int  <= 'h11c7; // Code pointer for 5_6
    9: romdata_int  <= 'h14b5; // Code pointer for 8_9
    10: romdata_int <= 'h1749; // Code pointer for 9_10
    11: romdata_int <= 'h19e3; // Code pointer for 1_5s
    12: romdata_int <= 'h1a2b; // Code pointer for 1_3s
    13: romdata_int <= 'h1a94; // Code pointer for 2_5s
    14: romdata_int <= 'h1b12; // Code pointer for 4_9s
    15: romdata_int <= 'h1b7b; // Code pointer for 3_5s
    16: romdata_int <= 'h1c38; // Code pointer for 2_3s
    17: romdata_int <= 'h1cce; // Code pointer for 11_15s
    18: romdata_int <= 'h1d5b; // Code pointer for 7_9s
    19: romdata_int <= 'h1de7; // Code pointer for 37_45s
    20: romdata_int <= 'h1e85; // Code pointer for 8_9s
    21: romdata_int <= 'h1687; // Line Descriptor
    22: romdata_int <= 'he8ae;
    23: romdata_int <= 'h6b0b;
    24: romdata_int <= 'h7808;
    25: romdata_int <= 'hd0d5;
    26: romdata_int <= 'h7486;
    27: romdata_int <= 'h1e89;
    28: romdata_int <= 'h202e;
    29: romdata_int <= 'h4;
    30: romdata_int <= 'h3b37;
    31: romdata_int <= 'hb29a;
    32: romdata_int <= 'h54b0;
    33: romdata_int <= 'hd95c;
    34: romdata_int <= 'h1687; // Line Descriptor
    35: romdata_int <= 'ha879;
    36: romdata_int <= 'hb0b8;
    37: romdata_int <= 'h87b;
    38: romdata_int <= 'hce7f;
    39: romdata_int <= 'h10a38;
    40: romdata_int <= 'h2cb9;
    41: romdata_int <= 'h7d3b;
    42: romdata_int <= 'hec7c;
    43: romdata_int <= 'hb702;
    44: romdata_int <= 'hea9b;
    45: romdata_int <= 'h4512;
    46: romdata_int <= 'h4a99;
    47: romdata_int <= 'h1687; // Line Descriptor
    48: romdata_int <= 'hee0d;
    49: romdata_int <= 'h10d28;
    50: romdata_int <= 'h948a;
    51: romdata_int <= 'h3a6b;
    52: romdata_int <= 'hc667;
    53: romdata_int <= 'h5855;
    54: romdata_int <= 'h1661;
    55: romdata_int <= 'h8ed5;
    56: romdata_int <= 'h771e;
    57: romdata_int <= 'hb0a5;
    58: romdata_int <= 'h1ee0;
    59: romdata_int <= 'h6ee6;
    60: romdata_int <= 'h1687; // Line Descriptor
    61: romdata_int <= 'he4a4;
    62: romdata_int <= 'h812c;
    63: romdata_int <= 'hc8a7;
    64: romdata_int <= 'hf4a6;
    65: romdata_int <= 'h762d;
    66: romdata_int <= 'h10643;
    67: romdata_int <= 'h4d28;
    68: romdata_int <= 'h108b0;
    69: romdata_int <= 'h3642;
    70: romdata_int <= 'ha673;
    71: romdata_int <= 'he47c;
    72: romdata_int <= 'hbce5;
    73: romdata_int <= 'h1687; // Line Descriptor
    74: romdata_int <= 'h903b;
    75: romdata_int <= 'h492b;
    76: romdata_int <= 'h6464;
    77: romdata_int <= 'hac90;
    78: romdata_int <= 'h6936;
    79: romdata_int <= 'h36d5;
    80: romdata_int <= 'h9462;
    81: romdata_int <= 'hfcf2;
    82: romdata_int <= 'hdab6;
    83: romdata_int <= 'hac9;
    84: romdata_int <= 'ha154;
    85: romdata_int <= 'h3e4a;
    86: romdata_int <= 'h1687; // Line Descriptor
    87: romdata_int <= 'h512c;
    88: romdata_int <= 'ha749;
    89: romdata_int <= 'hc67;
    90: romdata_int <= 'h32a6;
    91: romdata_int <= 'h3ef2;
    92: romdata_int <= 'h5a88;
    93: romdata_int <= 'hd127;
    94: romdata_int <= 'hcbd;
    95: romdata_int <= 'h9a5c;
    96: romdata_int <= 'h10648;
    97: romdata_int <= 'h9322;
    98: romdata_int <= 'h10101;
    99: romdata_int <= 'h1687; // Line Descriptor
    100: romdata_int <= 'he270;
    101: romdata_int <= 'hd94f;
    102: romdata_int <= 'h5c25;
    103: romdata_int <= 'h314d;
    104: romdata_int <= 'ha152;
    105: romdata_int <= 'h3d38;
    106: romdata_int <= 'hde8f;
    107: romdata_int <= 'h40e;
    108: romdata_int <= 'h48ab;
    109: romdata_int <= 'h8275;
    110: romdata_int <= 'h7241;
    111: romdata_int <= 'h604c;
    112: romdata_int <= 'h1687; // Line Descriptor
    113: romdata_int <= 'h924d;
    114: romdata_int <= 'h2148;
    115: romdata_int <= 'hca1a;
    116: romdata_int <= 'h1040a;
    117: romdata_int <= 'h6716;
    118: romdata_int <= 'hf8ee;
    119: romdata_int <= 'h5e66;
    120: romdata_int <= 'h10a32;
    121: romdata_int <= 'haef3;
    122: romdata_int <= 'h392a;
    123: romdata_int <= 'hc558;
    124: romdata_int <= 'h7858;
    125: romdata_int <= 'h1687; // Line Descriptor
    126: romdata_int <= 'hb431;
    127: romdata_int <= 'h44a0;
    128: romdata_int <= 'h8cd0;
    129: romdata_int <= 'h2344;
    130: romdata_int <= 'haa06;
    131: romdata_int <= 'h8630;
    132: romdata_int <= 'h5a9b;
    133: romdata_int <= 'h30d6;
    134: romdata_int <= 'h18df;
    135: romdata_int <= 'hacbe;
    136: romdata_int <= 'h2735;
    137: romdata_int <= 'h6854;
    138: romdata_int <= 'h1687; // Line Descriptor
    139: romdata_int <= 'h108a2;
    140: romdata_int <= 'h8a2a;
    141: romdata_int <= 'h96c9;
    142: romdata_int <= 'h24ce;
    143: romdata_int <= 'h4afd;
    144: romdata_int <= 'h7319;
    145: romdata_int <= 'he650;
    146: romdata_int <= 'he233;
    147: romdata_int <= 'h581c;
    148: romdata_int <= 'h1538;
    149: romdata_int <= 'h4e21;
    150: romdata_int <= 'hc708;
    151: romdata_int <= 'h1687; // Line Descriptor
    152: romdata_int <= 'h143f;
    153: romdata_int <= 'hde08;
    154: romdata_int <= 'he65;
    155: romdata_int <= 'h46e5;
    156: romdata_int <= 'h2ec0;
    157: romdata_int <= 'hec5d;
    158: romdata_int <= 'hf27b;
    159: romdata_int <= 'hd4fd;
    160: romdata_int <= 'hceeb;
    161: romdata_int <= 'hc818;
    162: romdata_int <= 'hd640;
    163: romdata_int <= 'h9722;
    164: romdata_int <= 'h1687; // Line Descriptor
    165: romdata_int <= 'h9e8c;
    166: romdata_int <= 'h607e;
    167: romdata_int <= 'h833f;
    168: romdata_int <= 'h7a1f;
    169: romdata_int <= 'h8823;
    170: romdata_int <= 'h2946;
    171: romdata_int <= 'h1c90;
    172: romdata_int <= 'ha2da;
    173: romdata_int <= 'h963;
    174: romdata_int <= 'h6c70;
    175: romdata_int <= 'h42b4;
    176: romdata_int <= 'h628f;
    177: romdata_int <= 'h1687; // Line Descriptor
    178: romdata_int <= 'hb27b;
    179: romdata_int <= 'h163e;
    180: romdata_int <= 'h9adb;
    181: romdata_int <= 'h9958;
    182: romdata_int <= 'hbcee;
    183: romdata_int <= 'h26c3;
    184: romdata_int <= 'hb445;
    185: romdata_int <= 'h8687;
    186: romdata_int <= 'h225c;
    187: romdata_int <= 'h5cca;
    188: romdata_int <= 'hc106;
    189: romdata_int <= 'hf37;
    190: romdata_int <= 'h1687; // Line Descriptor
    191: romdata_int <= 'hea73;
    192: romdata_int <= 'h842b;
    193: romdata_int <= 'h6358;
    194: romdata_int <= 'h100c5;
    195: romdata_int <= 'h52ad;
    196: romdata_int <= 'hcc35;
    197: romdata_int <= 'h8042;
    198: romdata_int <= 'h6617;
    199: romdata_int <= 'h3315;
    200: romdata_int <= 'h74c;
    201: romdata_int <= 'h6b06;
    202: romdata_int <= 'h5264;
    203: romdata_int <= 'h1687; // Line Descriptor
    204: romdata_int <= 'h7f3d;
    205: romdata_int <= 'h1aed;
    206: romdata_int <= 'hd731;
    207: romdata_int <= 'h391f;
    208: romdata_int <= 'hdcc4;
    209: romdata_int <= 'h414;
    210: romdata_int <= 'hfac9;
    211: romdata_int <= 'h1035b;
    212: romdata_int <= 'hee0a;
    213: romdata_int <= 'hc29a;
    214: romdata_int <= 'h2acb;
    215: romdata_int <= 'h9d1d;
    216: romdata_int <= 'h487; // Line Descriptor
    217: romdata_int <= 'h18a4;
    218: romdata_int <= 'hc0b3;
    219: romdata_int <= 'h7c3d;
    220: romdata_int <= 'h487; // Line Descriptor
    221: romdata_int <= 'h548f;
    222: romdata_int <= 'hf649;
    223: romdata_int <= 'hfecd;
    224: romdata_int <= 'h487; // Line Descriptor
    225: romdata_int <= 'h3503;
    226: romdata_int <= 'h122f;
    227: romdata_int <= 'ha2f8;
    228: romdata_int <= 'h487; // Line Descriptor
    229: romdata_int <= 'ha4dc;
    230: romdata_int <= 'hbee4;
    231: romdata_int <= 'hbada;
    232: romdata_int <= 'h487; // Line Descriptor
    233: romdata_int <= 'hc444;
    234: romdata_int <= 'h5f67;
    235: romdata_int <= 'h4e6a;
    236: romdata_int <= 'h487; // Line Descriptor
    237: romdata_int <= 'hfd19;
    238: romdata_int <= 'he61e;
    239: romdata_int <= 'h745;
    240: romdata_int <= 'h487; // Line Descriptor
    241: romdata_int <= 'h563f;
    242: romdata_int <= 'hc2f5;
    243: romdata_int <= 'hf0fe;
    244: romdata_int <= 'h487; // Line Descriptor
    245: romdata_int <= 'hfaa6;
    246: romdata_int <= 'h70d5;
    247: romdata_int <= 'h6eb1;
    248: romdata_int <= 'h487; // Line Descriptor
    249: romdata_int <= 'h6c97;
    250: romdata_int <= 'he01d;
    251: romdata_int <= 'h2ab3;
    252: romdata_int <= 'h487; // Line Descriptor
    253: romdata_int <= 'h111e;
    254: romdata_int <= 'hae3c;
    255: romdata_int <= 'h40e5;
    256: romdata_int <= 'h487; // Line Descriptor
    257: romdata_int <= 'h4307;
    258: romdata_int <= 'hb45;
    259: romdata_int <= 'h1029e;
    260: romdata_int <= 'h487; // Line Descriptor
    261: romdata_int <= 'h8e34;
    262: romdata_int <= 'hf351;
    263: romdata_int <= 'h9c6f;
    264: romdata_int <= 'h487; // Line Descriptor
    265: romdata_int <= 'hd228;
    266: romdata_int <= 'h45;
    267: romdata_int <= 'h4ca2;
    268: romdata_int <= 'h487; // Line Descriptor
    269: romdata_int <= 'h30b;
    270: romdata_int <= 'hdaf3;
    271: romdata_int <= 'hb657;
    272: romdata_int <= 'h487; // Line Descriptor
    273: romdata_int <= 'h1c36;
    274: romdata_int <= 'hb926;
    275: romdata_int <= 'hd4f9;
    276: romdata_int <= 'h487; // Line Descriptor
    277: romdata_int <= 'h3c7d;
    278: romdata_int <= 'hfedd;
    279: romdata_int <= 'h2860;
    280: romdata_int <= 'h487; // Line Descriptor
    281: romdata_int <= 'hca52;
    282: romdata_int <= 'ha8af;
    283: romdata_int <= 'h64a6;
    284: romdata_int <= 'h487; // Line Descriptor
    285: romdata_int <= 'he8ff;
    286: romdata_int <= 'ha449;
    287: romdata_int <= 'hab49;
    288: romdata_int <= 'h487; // Line Descriptor
    289: romdata_int <= 'h10467;
    290: romdata_int <= 'h855e;
    291: romdata_int <= 'h5041;
    292: romdata_int <= 'h487; // Line Descriptor
    293: romdata_int <= 'h906f;
    294: romdata_int <= 'hf550;
    295: romdata_int <= 'h34b5;
    296: romdata_int <= 'h487; // Line Descriptor
    297: romdata_int <= 'h10e2;
    298: romdata_int <= 'h2d11;
    299: romdata_int <= 'h8a06;
    300: romdata_int <= 'h487; // Line Descriptor
    301: romdata_int <= 'h2e38;
    302: romdata_int <= 'h10c62;
    303: romdata_int <= 'h40b4;
    304: romdata_int <= 'h487; // Line Descriptor
    305: romdata_int <= 'h5603;
    306: romdata_int <= 'h70c8;
    307: romdata_int <= 'hb822;
    308: romdata_int <= 'h487; // Line Descriptor
    309: romdata_int <= 'h8859;
    310: romdata_int <= 'h74e8;
    311: romdata_int <= 'h8ca0;
    312: romdata_int <= 'h487; // Line Descriptor
    313: romdata_int <= 'h9e08;
    314: romdata_int <= 'h9885;
    315: romdata_int <= 'h7a10;
    316: romdata_int <= 'h487; // Line Descriptor
    317: romdata_int <= 'h247e;
    318: romdata_int <= 'hd31e;
    319: romdata_int <= 'h4645;
    320: romdata_int <= 'h487; // Line Descriptor
    321: romdata_int <= 'h7e80;
    322: romdata_int <= 'hbeb5;
    323: romdata_int <= 'h12db;
    324: romdata_int <= 'h487; // Line Descriptor
    325: romdata_int <= 'hbb55;
    326: romdata_int <= 'hf8e5;
    327: romdata_int <= 'h1af3;
    328: romdata_int <= 'h487; // Line Descriptor
    329: romdata_int <= 'hf696;
    330: romdata_int <= 'he111;
    331: romdata_int <= 'hf087;
    332: romdata_int <= 'h587; // Line Descriptor
    333: romdata_int <= 'hdd59;
    334: romdata_int <= 'hcc98;
    335: romdata_int <= 'h2f3;
    336: romdata_int <= 'h1678; // Line Descriptor
    337: romdata_int <= 'hcf22;
    338: romdata_int <= 'h5eae;
    339: romdata_int <= 'h6b0b;
    340: romdata_int <= 'hb808;
    341: romdata_int <= 'h66d5;
    342: romdata_int <= 'h1a86;
    343: romdata_int <= 'h1c89;
    344: romdata_int <= 'h2e;
    345: romdata_int <= 'h3404;
    346: romdata_int <= 'h9f37;
    347: romdata_int <= 'h4c9a;
    348: romdata_int <= 'hb0;
    349: romdata_int <= 'h1678; // Line Descriptor
    350: romdata_int <= 'he860;
    351: romdata_int <= 'h9479;
    352: romdata_int <= 'h9cb8;
    353: romdata_int <= 'h67b;
    354: romdata_int <= 'hba7f;
    355: romdata_int <= 'hec38;
    356: romdata_int <= 'h2cb9;
    357: romdata_int <= 'h713b;
    358: romdata_int <= 'hd27c;
    359: romdata_int <= 'ha302;
    360: romdata_int <= 'hd09b;
    361: romdata_int <= 'h3d12;
    362: romdata_int <= 'h1678; // Line Descriptor
    363: romdata_int <= 'h6291;
    364: romdata_int <= 'hd20d;
    365: romdata_int <= 'hef28;
    366: romdata_int <= 'h808a;
    367: romdata_int <= 'h366b;
    368: romdata_int <= 'hb267;
    369: romdata_int <= 'h5255;
    370: romdata_int <= 'h1461;
    371: romdata_int <= 'h7cd5;
    372: romdata_int <= 'h691e;
    373: romdata_int <= 'h9ca5;
    374: romdata_int <= 'h1ce0;
    375: romdata_int <= 'h1678; // Line Descriptor
    376: romdata_int <= 'h96f3;
    377: romdata_int <= 'hc8a4;
    378: romdata_int <= 'h712c;
    379: romdata_int <= 'hb2a7;
    380: romdata_int <= 'hdaa6;
    381: romdata_int <= 'h722d;
    382: romdata_int <= 'hea43;
    383: romdata_int <= 'h4528;
    384: romdata_int <= 'heab0;
    385: romdata_int <= 'h2e42;
    386: romdata_int <= 'h9273;
    387: romdata_int <= 'hc87c;
    388: romdata_int <= 'h1678; // Line Descriptor
    389: romdata_int <= 'h9052;
    390: romdata_int <= 'h7e3b;
    391: romdata_int <= 'h3f2b;
    392: romdata_int <= 'h5664;
    393: romdata_int <= 'ha090;
    394: romdata_int <= 'h6b36;
    395: romdata_int <= 'h38d5;
    396: romdata_int <= 'h8662;
    397: romdata_int <= 'he0f2;
    398: romdata_int <= 'hc0b6;
    399: romdata_int <= 'hac9;
    400: romdata_int <= 'h8d54;
    401: romdata_int <= 'h1678; // Line Descriptor
    402: romdata_int <= 'h2b53;
    403: romdata_int <= 'h472c;
    404: romdata_int <= 'h9949;
    405: romdata_int <= 'hc67;
    406: romdata_int <= 'h34a6;
    407: romdata_int <= 'h40f2;
    408: romdata_int <= 'h5a88;
    409: romdata_int <= 'hbf27;
    410: romdata_int <= 'hcbd;
    411: romdata_int <= 'h845c;
    412: romdata_int <= 'he848;
    413: romdata_int <= 'h7f22;
    414: romdata_int <= 'h1678; // Line Descriptor
    415: romdata_int <= 'haa9f;
    416: romdata_int <= 'hcc82;
    417: romdata_int <= 'hc070;
    418: romdata_int <= 'h4d4f;
    419: romdata_int <= 'h3225;
    420: romdata_int <= 'h954d;
    421: romdata_int <= 'h3d52;
    422: romdata_int <= 'hc938;
    423: romdata_int <= 'h48f;
    424: romdata_int <= 'h400e;
    425: romdata_int <= 'h72ab;
    426: romdata_int <= 'hc475;
    427: romdata_int <= 'h1678; // Line Descriptor
    428: romdata_int <= 'h2505;
    429: romdata_int <= 'h2ca1;
    430: romdata_int <= 'h7a4d;
    431: romdata_int <= 'h1f48;
    432: romdata_int <= 'hb61a;
    433: romdata_int <= 'he80a;
    434: romdata_int <= 'h6316;
    435: romdata_int <= 'hdcee;
    436: romdata_int <= 'h5466;
    437: romdata_int <= 'hec32;
    438: romdata_int <= 'h98f3;
    439: romdata_int <= 'h372a;
    440: romdata_int <= 'h1678; // Line Descriptor
    441: romdata_int <= 'hd05f;
    442: romdata_int <= 'h34fe;
    443: romdata_int <= 'heca2;
    444: romdata_int <= 'h782a;
    445: romdata_int <= 'h88c9;
    446: romdata_int <= 'h24ce;
    447: romdata_int <= 'h4afd;
    448: romdata_int <= 'h6f19;
    449: romdata_int <= 'hc650;
    450: romdata_int <= 'hbe33;
    451: romdata_int <= 'h4a1c;
    452: romdata_int <= 'h1738;
    453: romdata_int <= 'h1678; // Line Descriptor
    454: romdata_int <= 'h1321;
    455: romdata_int <= 'hacc0;
    456: romdata_int <= 'h163f;
    457: romdata_int <= 'hc408;
    458: romdata_int <= 'he65;
    459: romdata_int <= 'h4ce5;
    460: romdata_int <= 'h30c0;
    461: romdata_int <= 'hd25d;
    462: romdata_int <= 'hd67b;
    463: romdata_int <= 'hb6fd;
    464: romdata_int <= 'hb2eb;
    465: romdata_int <= 'hac18;
    466: romdata_int <= 'h1678; // Line Descriptor
    467: romdata_int <= 'h2861;
    468: romdata_int <= 'hbc7f;
    469: romdata_int <= 'h868c;
    470: romdata_int <= 'h507e;
    471: romdata_int <= 'h7f3f;
    472: romdata_int <= 'h741f;
    473: romdata_int <= 'h8223;
    474: romdata_int <= 'h2746;
    475: romdata_int <= 'h1a90;
    476: romdata_int <= 'h8ada;
    477: romdata_int <= 'h963;
    478: romdata_int <= 'h5c70;
    479: romdata_int <= 'h1678; // Line Descriptor
    480: romdata_int <= 'h7306;
    481: romdata_int <= 'h5a0b;
    482: romdata_int <= 'h887b;
    483: romdata_int <= 'h1a3e;
    484: romdata_int <= 'h8cdb;
    485: romdata_int <= 'h8558;
    486: romdata_int <= 'ha6ee;
    487: romdata_int <= 'h2ac3;
    488: romdata_int <= 'h9445;
    489: romdata_int <= 'h6e87;
    490: romdata_int <= 'h1e5c;
    491: romdata_int <= 'h4eca;
    492: romdata_int <= 'h1678; // Line Descriptor
    493: romdata_int <= 'hae82;
    494: romdata_int <= 'hd667;
    495: romdata_int <= 'hd473;
    496: romdata_int <= 'h6e2b;
    497: romdata_int <= 'h6158;
    498: romdata_int <= 'he6c5;
    499: romdata_int <= 'h50ad;
    500: romdata_int <= 'hae35;
    501: romdata_int <= 'h6442;
    502: romdata_int <= 'h5617;
    503: romdata_int <= 'h2d15;
    504: romdata_int <= 'h74c;
    505: romdata_int <= 'h1678; // Line Descriptor
    506: romdata_int <= 'ha62c;
    507: romdata_int <= 'h3abb;
    508: romdata_int <= 'h673d;
    509: romdata_int <= 'h22ed;
    510: romdata_int <= 'hc131;
    511: romdata_int <= 'h3f1f;
    512: romdata_int <= 'hc6c4;
    513: romdata_int <= 'h814;
    514: romdata_int <= 'hdac9;
    515: romdata_int <= 'he55b;
    516: romdata_int <= 'hc20a;
    517: romdata_int <= 'ha69a;
    518: romdata_int <= 'h1678; // Line Descriptor
    519: romdata_int <= 'h921e;
    520: romdata_int <= 'h8d45;
    521: romdata_int <= 'ha078;
    522: romdata_int <= 'h4efc;
    523: romdata_int <= 'h5738;
    524: romdata_int <= 'h283f;
    525: romdata_int <= 'heef5;
    526: romdata_int <= 'h4efe;
    527: romdata_int <= 'hdf4b;
    528: romdata_int <= 'hb8a8;
    529: romdata_int <= 'h1897;
    530: romdata_int <= 'hb4a6;
    531: romdata_int <= 'h1678; // Line Descriptor
    532: romdata_int <= 'h851e;
    533: romdata_int <= 'h683c;
    534: romdata_int <= 'h5ce5;
    535: romdata_int <= 'hdc6b;
    536: romdata_int <= 'h4639;
    537: romdata_int <= 'h7966;
    538: romdata_int <= 'hd07;
    539: romdata_int <= 'h8b45;
    540: romdata_int <= 'h329e;
    541: romdata_int <= 'h7a81;
    542: romdata_int <= 'h794d;
    543: romdata_int <= 'h468b;
    544: romdata_int <= 'h1678; // Line Descriptor
    545: romdata_int <= 'h520e;
    546: romdata_int <= 'h1937;
    547: romdata_int <= 'he34c;
    548: romdata_int <= 'h3c91;
    549: romdata_int <= 'hbd0b;
    550: romdata_int <= 'h4f3;
    551: romdata_int <= 'h6457;
    552: romdata_int <= 'h166c;
    553: romdata_int <= 'h2aee;
    554: romdata_int <= 'h66f4;
    555: romdata_int <= 'h1236;
    556: romdata_int <= 'hcf26;
    557: romdata_int <= 'h1678; // Line Descriptor
    558: romdata_int <= 'h2006;
    559: romdata_int <= 'h7c3a;
    560: romdata_int <= 'hdb60;
    561: romdata_int <= 'h2e49;
    562: romdata_int <= 'h5e38;
    563: romdata_int <= 'hde62;
    564: romdata_int <= 'h96b4;
    565: romdata_int <= 'ha56;
    566: romdata_int <= 'h3860;
    567: romdata_int <= 'h74d8;
    568: romdata_int <= 'h8e03;
    569: romdata_int <= 'haac8;
    570: romdata_int <= 'h1678; // Line Descriptor
    571: romdata_int <= 'ha10;
    572: romdata_int <= 'h5458;
    573: romdata_int <= 'h32ee;
    574: romdata_int <= 'h6465;
    575: romdata_int <= 'h487e;
    576: romdata_int <= 'ha91e;
    577: romdata_int <= 'h8e45;
    578: romdata_int <= 'h926e;
    579: romdata_int <= 'h60a8;
    580: romdata_int <= 'h5030;
    581: romdata_int <= 'he80;
    582: romdata_int <= 'h58b5;
    583: romdata_int <= 'h1678; // Line Descriptor
    584: romdata_int <= 'h9e87;
    585: romdata_int <= 'h413b;
    586: romdata_int <= 'he121;
    587: romdata_int <= 'h14b1;
    588: romdata_int <= 'he11c;
    589: romdata_int <= 'hac3d;
    590: romdata_int <= 'hb159;
    591: romdata_int <= 'hd498;
    592: romdata_int <= 'h86f3;
    593: romdata_int <= 'haed9;
    594: romdata_int <= 'h6ad4;
    595: romdata_int <= 'hb03a;
    596: romdata_int <= 'h478; // Line Descriptor
    597: romdata_int <= 'hd94c;
    598: romdata_int <= 'h3aeb;
    599: romdata_int <= 'h76cf;
    600: romdata_int <= 'h478; // Line Descriptor
    601: romdata_int <= 'h1091;
    602: romdata_int <= 'he476;
    603: romdata_int <= 'he344;
    604: romdata_int <= 'h478; // Line Descriptor
    605: romdata_int <= 'h1d43;
    606: romdata_int <= 'h1085;
    607: romdata_int <= 'h26ed;
    608: romdata_int <= 'h478; // Line Descriptor
    609: romdata_int <= 'h959;
    610: romdata_int <= 'h12e3;
    611: romdata_int <= 'h82e4;
    612: romdata_int <= 'h478; // Line Descriptor
    613: romdata_int <= 'h8b57;
    614: romdata_int <= 'ha432;
    615: romdata_int <= 'h4567;
    616: romdata_int <= 'h478; // Line Descriptor
    617: romdata_int <= 'h4a74;
    618: romdata_int <= 'h7629;
    619: romdata_int <= 'hbd52;
    620: romdata_int <= 'h478; // Line Descriptor
    621: romdata_int <= 'hba19;
    622: romdata_int <= 'h9c1c;
    623: romdata_int <= 'h9123;
    624: romdata_int <= 'h478; // Line Descriptor
    625: romdata_int <= 'h51c;
    626: romdata_int <= 'h6833;
    627: romdata_int <= 'ha0ef;
    628: romdata_int <= 'h478; // Line Descriptor
    629: romdata_int <= 'hb55f;
    630: romdata_int <= 'h7b1c;
    631: romdata_int <= 'hcb55;
    632: romdata_int <= 'h478; // Line Descriptor
    633: romdata_int <= 'h827a;
    634: romdata_int <= 'h2e94;
    635: romdata_int <= 'h6c54;
    636: romdata_int <= 'h478; // Line Descriptor
    637: romdata_int <= 'he75b;
    638: romdata_int <= 'h594c;
    639: romdata_int <= 'hbabd;
    640: romdata_int <= 'h478; // Line Descriptor
    641: romdata_int <= 'hbe79;
    642: romdata_int <= 'he281;
    643: romdata_int <= 'ha40d;
    644: romdata_int <= 'h478; // Line Descriptor
    645: romdata_int <= 'h8ef2;
    646: romdata_int <= 'hcb34;
    647: romdata_int <= 'h294c;
    648: romdata_int <= 'h478; // Line Descriptor
    649: romdata_int <= 'hc64f;
    650: romdata_int <= 'h9117;
    651: romdata_int <= 'h4205;
    652: romdata_int <= 'h478; // Line Descriptor
    653: romdata_int <= 'hde6b;
    654: romdata_int <= 'h22b0;
    655: romdata_int <= 'h114a;
    656: romdata_int <= 'h478; // Line Descriptor
    657: romdata_int <= 'ha93e;
    658: romdata_int <= 'h2e4;
    659: romdata_int <= 'h22f5;
    660: romdata_int <= 'h478; // Line Descriptor
    661: romdata_int <= 'h7618;
    662: romdata_int <= 'hb854;
    663: romdata_int <= 'hef2f;
    664: romdata_int <= 'h478; // Line Descriptor
    665: romdata_int <= 'h6cf2;
    666: romdata_int <= 'h9a2c;
    667: romdata_int <= 'h30a0;
    668: romdata_int <= 'h478; // Line Descriptor
    669: romdata_int <= 'ha44f;
    670: romdata_int <= 'h98cb;
    671: romdata_int <= 'h9aee;
    672: romdata_int <= 'h478; // Line Descriptor
    673: romdata_int <= 'hc34e;
    674: romdata_int <= 'h5c13;
    675: romdata_int <= 'h8070;
    676: romdata_int <= 'h478; // Line Descriptor
    677: romdata_int <= 'he438;
    678: romdata_int <= 'hceb3;
    679: romdata_int <= 'h4962;
    680: romdata_int <= 'h478; // Line Descriptor
    681: romdata_int <= 'hb752;
    682: romdata_int <= 'hb564;
    683: romdata_int <= 'h3ad6;
    684: romdata_int <= 'h478; // Line Descriptor
    685: romdata_int <= 'heb06;
    686: romdata_int <= 'hc50b;
    687: romdata_int <= 'hcd3d;
    688: romdata_int <= 'h478; // Line Descriptor
    689: romdata_int <= 'h309b;
    690: romdata_int <= 'hd75c;
    691: romdata_int <= 'h7147;
    692: romdata_int <= 'h478; // Line Descriptor
    693: romdata_int <= 'h139;
    694: romdata_int <= 'h1e77;
    695: romdata_int <= 'h5a87;
    696: romdata_int <= 'h478; // Line Descriptor
    697: romdata_int <= 'hca38;
    698: romdata_int <= 'h9eb4;
    699: romdata_int <= 'h1507;
    700: romdata_int <= 'h478; // Line Descriptor
    701: romdata_int <= 'h26d3;
    702: romdata_int <= 'h6d1;
    703: romdata_int <= 'h2b8;
    704: romdata_int <= 'h478; // Line Descriptor
    705: romdata_int <= 'he43;
    706: romdata_int <= 'hc205;
    707: romdata_int <= 'hd925;
    708: romdata_int <= 'h478; // Line Descriptor
    709: romdata_int <= 'h5852;
    710: romdata_int <= 'h428e;
    711: romdata_int <= 'h96a6;
    712: romdata_int <= 'h478; // Line Descriptor
    713: romdata_int <= 'hb0df;
    714: romdata_int <= 'hab25;
    715: romdata_int <= 'hdc45;
    716: romdata_int <= 'h478; // Line Descriptor
    717: romdata_int <= 'h749b;
    718: romdata_int <= 'h6c86;
    719: romdata_int <= 'h5e7b;
    720: romdata_int <= 'h478; // Line Descriptor
    721: romdata_int <= 'ha265;
    722: romdata_int <= 'h8112;
    723: romdata_int <= 'he629;
    724: romdata_int <= 'h478; // Line Descriptor
    725: romdata_int <= 'h48d2;
    726: romdata_int <= 'h200a;
    727: romdata_int <= 'hd544;
    728: romdata_int <= 'h478; // Line Descriptor
    729: romdata_int <= 'h4566;
    730: romdata_int <= 'h7cce;
    731: romdata_int <= 'h5248;
    732: romdata_int <= 'h478; // Line Descriptor
    733: romdata_int <= 'h2ec;
    734: romdata_int <= 'h1829;
    735: romdata_int <= 'h631d;
    736: romdata_int <= 'h478; // Line Descriptor
    737: romdata_int <= 'h3622;
    738: romdata_int <= 'hccf4;
    739: romdata_int <= 'ha90b;
    740: romdata_int <= 'h478; // Line Descriptor
    741: romdata_int <= 'h9ab8;
    742: romdata_int <= 'hd015;
    743: romdata_int <= 'h8878;
    744: romdata_int <= 'h478; // Line Descriptor
    745: romdata_int <= 'h3943;
    746: romdata_int <= 'ha2e1;
    747: romdata_int <= 'h2042;
    748: romdata_int <= 'h478; // Line Descriptor
    749: romdata_int <= 'h6024;
    750: romdata_int <= 'hd8d9;
    751: romdata_int <= 'h2458;
    752: romdata_int <= 'h578; // Line Descriptor
    753: romdata_int <= 'h42d3;
    754: romdata_int <= 'h5422;
    755: romdata_int <= 'h3f4b;
    756: romdata_int <= 'h166c; // Line Descriptor
    757: romdata_int <= 'hbb22;
    758: romdata_int <= 'h54ae;
    759: romdata_int <= 'h610b;
    760: romdata_int <= 'ha608;
    761: romdata_int <= 'h5cd5;
    762: romdata_int <= 'h1886;
    763: romdata_int <= 'h1a89;
    764: romdata_int <= 'h2e;
    765: romdata_int <= 'h2e04;
    766: romdata_int <= 'h8f37;
    767: romdata_int <= 'h449a;
    768: romdata_int <= 'hb0;
    769: romdata_int <= 'h166c; // Line Descriptor
    770: romdata_int <= 'hd079;
    771: romdata_int <= 'h86b8;
    772: romdata_int <= 'h8c7b;
    773: romdata_int <= 'h67f;
    774: romdata_int <= 'ha838;
    775: romdata_int <= 'hd4b9;
    776: romdata_int <= 'h293b;
    777: romdata_int <= 'h647c;
    778: romdata_int <= 'hbd02;
    779: romdata_int <= 'h929b;
    780: romdata_int <= 'h3712;
    781: romdata_int <= 'h3a99;
    782: romdata_int <= 'h166c; // Line Descriptor
    783: romdata_int <= 'hbe0d;
    784: romdata_int <= 'hd728;
    785: romdata_int <= 'h748a;
    786: romdata_int <= 'h2c6b;
    787: romdata_int <= 'ha067;
    788: romdata_int <= 'h4a55;
    789: romdata_int <= 'h1261;
    790: romdata_int <= 'h74d5;
    791: romdata_int <= 'h611e;
    792: romdata_int <= 'h90a5;
    793: romdata_int <= 'h18e0;
    794: romdata_int <= 'h5ae6;
    795: romdata_int <= 'h166c; // Line Descriptor
    796: romdata_int <= 'hb52c;
    797: romdata_int <= 'h64a7;
    798: romdata_int <= 'h9ea6;
    799: romdata_int <= 'hc22d;
    800: romdata_int <= 'h6243;
    801: romdata_int <= 'hd328;
    802: romdata_int <= 'h3cb0;
    803: romdata_int <= 'h3042;
    804: romdata_int <= 'h8473;
    805: romdata_int <= 'hb67c;
    806: romdata_int <= 'h98e5;
    807: romdata_int <= 'h66c9;
    808: romdata_int <= 'h166c; // Line Descriptor
    809: romdata_int <= 'h3b2b;
    810: romdata_int <= 'h4e64;
    811: romdata_int <= 'h8890;
    812: romdata_int <= 'h5336;
    813: romdata_int <= 'h34d5;
    814: romdata_int <= 'h7c62;
    815: romdata_int <= 'hc8f2;
    816: romdata_int <= 'hb0b6;
    817: romdata_int <= 'hac9;
    818: romdata_int <= 'h8154;
    819: romdata_int <= 'h304a;
    820: romdata_int <= 'h2277;
    821: romdata_int <= 'h166c; // Line Descriptor
    822: romdata_int <= 'h8349;
    823: romdata_int <= 'ha67;
    824: romdata_int <= 'h28a6;
    825: romdata_int <= 'h30f2;
    826: romdata_int <= 'h5288;
    827: romdata_int <= 'ha727;
    828: romdata_int <= 'h8bd;
    829: romdata_int <= 'h805c;
    830: romdata_int <= 'hd448;
    831: romdata_int <= 'h7922;
    832: romdata_int <= 'hcd01;
    833: romdata_int <= 'hb934;
    834: romdata_int <= 'h166c; // Line Descriptor
    835: romdata_int <= 'haa82;
    836: romdata_int <= 'h4670;
    837: romdata_int <= 'h274f;
    838: romdata_int <= 'h7c25;
    839: romdata_int <= 'h394d;
    840: romdata_int <= 'hb552;
    841: romdata_int <= 'h538;
    842: romdata_int <= 'h3e8f;
    843: romdata_int <= 'h6c0e;
    844: romdata_int <= 'h3cab;
    845: romdata_int <= 'hb275;
    846: romdata_int <= 'h5e41;
    847: romdata_int <= 'h166c; // Line Descriptor
    848: romdata_int <= 'h24a1;
    849: romdata_int <= 'h704d;
    850: romdata_int <= 'h1b48;
    851: romdata_int <= 'ha01a;
    852: romdata_int <= 'hd00a;
    853: romdata_int <= 'h5916;
    854: romdata_int <= 'hc4ee;
    855: romdata_int <= 'h5066;
    856: romdata_int <= 'hd632;
    857: romdata_int <= 'h8af3;
    858: romdata_int <= 'h2b2a;
    859: romdata_int <= 'ha158;
    860: romdata_int <= 'h166c; // Line Descriptor
    861: romdata_int <= 'h348d;
    862: romdata_int <= 'h9231;
    863: romdata_int <= 'h38a0;
    864: romdata_int <= 'h6ed0;
    865: romdata_int <= 'h2344;
    866: romdata_int <= 'h8c06;
    867: romdata_int <= 'h7030;
    868: romdata_int <= 'h4c9b;
    869: romdata_int <= 'h26d6;
    870: romdata_int <= 'h10df;
    871: romdata_int <= 'h86be;
    872: romdata_int <= 'h1b35;
    873: romdata_int <= 'h166c; // Line Descriptor
    874: romdata_int <= 'h2efe;
    875: romdata_int <= 'hd4a2;
    876: romdata_int <= 'h6c2a;
    877: romdata_int <= 'h76c9;
    878: romdata_int <= 'h24ce;
    879: romdata_int <= 'h42fd;
    880: romdata_int <= 'h6919;
    881: romdata_int <= 'hb850;
    882: romdata_int <= 'hb033;
    883: romdata_int <= 'h481c;
    884: romdata_int <= 'hf38;
    885: romdata_int <= 'h4021;
    886: romdata_int <= 'h166c; // Line Descriptor
    887: romdata_int <= 'h9c3f;
    888: romdata_int <= 'h1208;
    889: romdata_int <= 'hb265;
    890: romdata_int <= 'hce5;
    891: romdata_int <= 'h44c0;
    892: romdata_int <= 'h2e5d;
    893: romdata_int <= 'hbe7b;
    894: romdata_int <= 'haafd;
    895: romdata_int <= 'ha6eb;
    896: romdata_int <= 'ha218;
    897: romdata_int <= 'hac40;
    898: romdata_int <= 'h7522;
    899: romdata_int <= 'h166c; // Line Descriptor
    900: romdata_int <= 'h7a8c;
    901: romdata_int <= 'h4a7e;
    902: romdata_int <= 'h633f;
    903: romdata_int <= 'h5a1f;
    904: romdata_int <= 'h7823;
    905: romdata_int <= 'h2746;
    906: romdata_int <= 'h1490;
    907: romdata_int <= 'h8eda;
    908: romdata_int <= 'h563;
    909: romdata_int <= 'h5670;
    910: romdata_int <= 'h3eb4;
    911: romdata_int <= 'h4e8f;
    912: romdata_int <= 'h166c; // Line Descriptor
    913: romdata_int <= 'h847b;
    914: romdata_int <= 'h163e;
    915: romdata_int <= 'h72db;
    916: romdata_int <= 'h6958;
    917: romdata_int <= 'h94ee;
    918: romdata_int <= 'h2cc3;
    919: romdata_int <= 'h7645;
    920: romdata_int <= 'h1087;
    921: romdata_int <= 'h945c;
    922: romdata_int <= 'h4cca;
    923: romdata_int <= 'h9f06;
    924: romdata_int <= 'h737;
    925: romdata_int <= 'h166c; // Line Descriptor
    926: romdata_int <= 'hbc73;
    927: romdata_int <= 'h662b;
    928: romdata_int <= 'h4d58;
    929: romdata_int <= 'hcec5;
    930: romdata_int <= 'h4ead;
    931: romdata_int <= 'h9c35;
    932: romdata_int <= 'h6c42;
    933: romdata_int <= 'h5a17;
    934: romdata_int <= 'h2915;
    935: romdata_int <= 'h94c;
    936: romdata_int <= 'h5506;
    937: romdata_int <= 'h4664;
    938: romdata_int <= 'h166c; // Line Descriptor
    939: romdata_int <= 'h5f3d;
    940: romdata_int <= 'h1ced;
    941: romdata_int <= 'had31;
    942: romdata_int <= 'h2b1f;
    943: romdata_int <= 'hb6c4;
    944: romdata_int <= 'ha14;
    945: romdata_int <= 'hc6c9;
    946: romdata_int <= 'hcd5b;
    947: romdata_int <= 'hbe0a;
    948: romdata_int <= 'h9c9a;
    949: romdata_int <= 'h1ecb;
    950: romdata_int <= 'h7b1d;
    951: romdata_int <= 'h166c; // Line Descriptor
    952: romdata_int <= 'h98fc;
    953: romdata_int <= 'h4538;
    954: romdata_int <= 'h403f;
    955: romdata_int <= 'h20f5;
    956: romdata_int <= 'hd6fe;
    957: romdata_int <= 'h494b;
    958: romdata_int <= 'hcaa8;
    959: romdata_int <= 'hac97;
    960: romdata_int <= 'h16a6;
    961: romdata_int <= 'hb4d5;
    962: romdata_int <= 'hc8b1;
    963: romdata_int <= 'h58a1;
    964: romdata_int <= 'h166c; // Line Descriptor
    965: romdata_int <= 'hc66b;
    966: romdata_int <= 'h3639;
    967: romdata_int <= 'h5966;
    968: romdata_int <= 'h907;
    969: romdata_int <= 'h7345;
    970: romdata_int <= 'h329e;
    971: romdata_int <= 'h8481;
    972: romdata_int <= 'h834d;
    973: romdata_int <= 'h508b;
    974: romdata_int <= 'hba99;
    975: romdata_int <= 'h2c34;
    976: romdata_int <= 'h8951;
    977: romdata_int <= 'h166c; // Line Descriptor
    978: romdata_int <= 'h4291;
    979: romdata_int <= 'haf0b;
    980: romdata_int <= 'h2f3;
    981: romdata_int <= 'h4857;
    982: romdata_int <= 'h166c;
    983: romdata_int <= 'h20ee;
    984: romdata_int <= 'h6af4;
    985: romdata_int <= 'hc36;
    986: romdata_int <= 'hc726;
    987: romdata_int <= 'hcf9;
    988: romdata_int <= 'hc44a;
    989: romdata_int <= 'hcb56;
    990: romdata_int <= 'h166c; // Line Descriptor
    991: romdata_int <= 'h14e2;
    992: romdata_int <= 'h56ff;
    993: romdata_int <= 'h9649;
    994: romdata_int <= 'h3d49;
    995: romdata_int <= 'h9f5d;
    996: romdata_int <= 'h90a4;
    997: romdata_int <= 'h5469;
    998: romdata_int <= 'h4067;
    999: romdata_int <= 'h6f5e;
    1000: romdata_int <= 'h6a41;
    1001: romdata_int <= 'haac8;
    1002: romdata_int <= 'h7f3f;
    1003: romdata_int <= 'h166c; // Line Descriptor
    1004: romdata_int <= 'h8a65;
    1005: romdata_int <= 'h327e;
    1006: romdata_int <= 'ha31e;
    1007: romdata_int <= 'h8045;
    1008: romdata_int <= 'h7e6e;
    1009: romdata_int <= 'h6ea8;
    1010: romdata_int <= 'h5e30;
    1011: romdata_int <= 'h280;
    1012: romdata_int <= 'h52b5;
    1013: romdata_int <= 'h12db;
    1014: romdata_int <= 'h3467;
    1015: romdata_int <= 'h8d49;
    1016: romdata_int <= 'h166c; // Line Descriptor
    1017: romdata_int <= 'h10b1;
    1018: romdata_int <= 'hcd1c;
    1019: romdata_int <= 'ha43d;
    1020: romdata_int <= 'ha959;
    1021: romdata_int <= 'hbc98;
    1022: romdata_int <= 'h92f3;
    1023: romdata_int <= 'ha4d9;
    1024: romdata_int <= 'h7ad4;
    1025: romdata_int <= 'ha83a;
    1026: romdata_int <= 'h633b;
    1027: romdata_int <= 'hc251;
    1028: romdata_int <= 'haeba;
    1029: romdata_int <= 'h166c; // Line Descriptor
    1030: romdata_int <= 'hcb43;
    1031: romdata_int <= 'h9a85;
    1032: romdata_int <= 'h90ed;
    1033: romdata_int <= 'h1826;
    1034: romdata_int <= 'hce1b;
    1035: romdata_int <= 'hc2c2;
    1036: romdata_int <= 'h6159;
    1037: romdata_int <= 'h46e3;
    1038: romdata_int <= 'hcee4;
    1039: romdata_int <= 'h20ba;
    1040: romdata_int <= 'h14e6;
    1041: romdata_int <= 'h2470;
    1042: romdata_int <= 'h166c; // Line Descriptor
    1043: romdata_int <= 'h7f61;
    1044: romdata_int <= 'h1f08;
    1045: romdata_int <= 'h5079;
    1046: romdata_int <= 'h6a81;
    1047: romdata_int <= 'h2a0d;
    1048: romdata_int <= 'hbac6;
    1049: romdata_int <= 'h371d;
    1050: romdata_int <= 'ha24f;
    1051: romdata_int <= 'hd2f2;
    1052: romdata_int <= 'hd134;
    1053: romdata_int <= 'h734c;
    1054: romdata_int <= 'h9b2c;
    1055: romdata_int <= 'h166c; // Line Descriptor
    1056: romdata_int <= 'h8e36;
    1057: romdata_int <= 'h5d3e;
    1058: romdata_int <= 'h22e4;
    1059: romdata_int <= 'hc0f5;
    1060: romdata_int <= 'h6d5;
    1061: romdata_int <= 'hb2fc;
    1062: romdata_int <= 'h1f62;
    1063: romdata_int <= 'h3a18;
    1064: romdata_int <= 'h6454;
    1065: romdata_int <= 'ha52f;
    1066: romdata_int <= 'h7cc7;
    1067: romdata_int <= 'h2ad;
    1068: romdata_int <= 'h46c; // Line Descriptor
    1069: romdata_int <= 'hea0;
    1070: romdata_int <= 'h98fc;
    1071: romdata_int <= 'h32b0;
    1072: romdata_int <= 'h46c; // Line Descriptor
    1073: romdata_int <= 'hb8ee;
    1074: romdata_int <= 'h5726;
    1075: romdata_int <= 'h7070;
    1076: romdata_int <= 'h46c; // Line Descriptor
    1077: romdata_int <= 'hb070;
    1078: romdata_int <= 'hc144;
    1079: romdata_int <= 'h1d21;
    1080: romdata_int <= 'h46c; // Line Descriptor
    1081: romdata_int <= 'h3f62;
    1082: romdata_int <= 'h1d35;
    1083: romdata_int <= 'h68e6;
    1084: romdata_int <= 'h46c; // Line Descriptor
    1085: romdata_int <= 'h4d6;
    1086: romdata_int <= 'haf5f;
    1087: romdata_int <= 'hc113;
    1088: romdata_int <= 'h46c; // Line Descriptor
    1089: romdata_int <= 'hc93d;
    1090: romdata_int <= 'h9661;
    1091: romdata_int <= 'h834f;
    1092: romdata_int <= 'h46c; // Line Descriptor
    1093: romdata_int <= 'hb747;
    1094: romdata_int <= 'h8601;
    1095: romdata_int <= 'h9642;
    1096: romdata_int <= 'h46c; // Line Descriptor
    1097: romdata_int <= 'h9487;
    1098: romdata_int <= 'h9b61;
    1099: romdata_int <= 'h42d1;
    1100: romdata_int <= 'h46c; // Line Descriptor
    1101: romdata_int <= 'h107;
    1102: romdata_int <= 'he3d;
    1103: romdata_int <= 'h5c09;
    1104: romdata_int <= 'h46c; // Line Descriptor
    1105: romdata_int <= 'h78b8;
    1106: romdata_int <= 'h8820;
    1107: romdata_int <= 'h4b0f;
    1108: romdata_int <= 'h46c; // Line Descriptor
    1109: romdata_int <= 'hd325;
    1110: romdata_int <= 'h66bb;
    1111: romdata_int <= 'h384b;
    1112: romdata_int <= 'h46c; // Line Descriptor
    1113: romdata_int <= 'hc4a6;
    1114: romdata_int <= 'h8b50;
    1115: romdata_int <= 'h76f7;
    1116: romdata_int <= 'h46c; // Line Descriptor
    1117: romdata_int <= 'hb645;
    1118: romdata_int <= 'h8713;
    1119: romdata_int <= 'hb07d;
    1120: romdata_int <= 'h46c; // Line Descriptor
    1121: romdata_int <= 'h627b;
    1122: romdata_int <= 'h5af0;
    1123: romdata_int <= 'h4e4e;
    1124: romdata_int <= 'h46c; // Line Descriptor
    1125: romdata_int <= 'h4086;
    1126: romdata_int <= 'h9954;
    1127: romdata_int <= 'h6cb6;
    1128: romdata_int <= 'h46c; // Line Descriptor
    1129: romdata_int <= 'hc829;
    1130: romdata_int <= 'h36ea;
    1131: romdata_int <= 'ha443;
    1132: romdata_int <= 'h46c; // Line Descriptor
    1133: romdata_int <= 'hc744;
    1134: romdata_int <= 'h7cec;
    1135: romdata_int <= 'h489;
    1136: romdata_int <= 'h46c; // Line Descriptor
    1137: romdata_int <= 'h6048;
    1138: romdata_int <= 'hd601;
    1139: romdata_int <= 'h780b;
    1140: romdata_int <= 'h46c; // Line Descriptor
    1141: romdata_int <= 'h891d;
    1142: romdata_int <= 'h8c31;
    1143: romdata_int <= 'h16a0;
    1144: romdata_int <= 'h46c; // Line Descriptor
    1145: romdata_int <= 'hc10b;
    1146: romdata_int <= 'h1318;
    1147: romdata_int <= 'h92fa;
    1148: romdata_int <= 'h46c; // Line Descriptor
    1149: romdata_int <= 'hcc78;
    1150: romdata_int <= 'h6613;
    1151: romdata_int <= 'hc96;
    1152: romdata_int <= 'h46c; // Line Descriptor
    1153: romdata_int <= 'h242;
    1154: romdata_int <= 'hbd28;
    1155: romdata_int <= 'h80b5;
    1156: romdata_int <= 'h46c; // Line Descriptor
    1157: romdata_int <= 'h1058;
    1158: romdata_int <= 'h18cb;
    1159: romdata_int <= 'h7b67;
    1160: romdata_int <= 'h46c; // Line Descriptor
    1161: romdata_int <= 'hcb4b;
    1162: romdata_int <= 'h7538;
    1163: romdata_int <= 'h1cd9;
    1164: romdata_int <= 'h46c; // Line Descriptor
    1165: romdata_int <= 'h2aad;
    1166: romdata_int <= 'h4909;
    1167: romdata_int <= 'h96a7;
    1168: romdata_int <= 'h46c; // Line Descriptor
    1169: romdata_int <= 'h8ad2;
    1170: romdata_int <= 'h30fe;
    1171: romdata_int <= 'h72a;
    1172: romdata_int <= 'h46c; // Line Descriptor
    1173: romdata_int <= 'h5305;
    1174: romdata_int <= 'h5125;
    1175: romdata_int <= 'h3917;
    1176: romdata_int <= 'h46c; // Line Descriptor
    1177: romdata_int <= 'h828d;
    1178: romdata_int <= 'h764e;
    1179: romdata_int <= 'h3d03;
    1180: romdata_int <= 'h46c; // Line Descriptor
    1181: romdata_int <= 'ha889;
    1182: romdata_int <= 'h647b;
    1183: romdata_int <= 'h7074;
    1184: romdata_int <= 'h46c; // Line Descriptor
    1185: romdata_int <= 'h3509;
    1186: romdata_int <= 'h9417;
    1187: romdata_int <= 'h3eb6;
    1188: romdata_int <= 'h46c; // Line Descriptor
    1189: romdata_int <= 'hce39;
    1190: romdata_int <= 'h8e29;
    1191: romdata_int <= 'hb8f3;
    1192: romdata_int <= 'h46c; // Line Descriptor
    1193: romdata_int <= 'h906e;
    1194: romdata_int <= 'hb506;
    1195: romdata_int <= 'hb24d;
    1196: romdata_int <= 'h46c; // Line Descriptor
    1197: romdata_int <= 'h3262;
    1198: romdata_int <= 'hc208;
    1199: romdata_int <= 'h2c46;
    1200: romdata_int <= 'h46c; // Line Descriptor
    1201: romdata_int <= 'h6e60;
    1202: romdata_int <= 'h1e7a;
    1203: romdata_int <= 'h44f8;
    1204: romdata_int <= 'h46c; // Line Descriptor
    1205: romdata_int <= 'h5c93;
    1206: romdata_int <= 'h5553;
    1207: romdata_int <= 'h84c6;
    1208: romdata_int <= 'h46c; // Line Descriptor
    1209: romdata_int <= 'h2061;
    1210: romdata_int <= 'h280e;
    1211: romdata_int <= 'h220b;
    1212: romdata_int <= 'h46c; // Line Descriptor
    1213: romdata_int <= 'hbf1a;
    1214: romdata_int <= 'had51;
    1215: romdata_int <= 'h1acd;
    1216: romdata_int <= 'h46c; // Line Descriptor
    1217: romdata_int <= 'ha02f;
    1218: romdata_int <= 'hc468;
    1219: romdata_int <= 'hf3d;
    1220: romdata_int <= 'h46c; // Line Descriptor
    1221: romdata_int <= 'hd108;
    1222: romdata_int <= 'h6b47;
    1223: romdata_int <= 'h4c7b;
    1224: romdata_int <= 'h46c; // Line Descriptor
    1225: romdata_int <= 'hd452;
    1226: romdata_int <= 'ha20d;
    1227: romdata_int <= 'h24c4;
    1228: romdata_int <= 'h46c; // Line Descriptor
    1229: romdata_int <= 'hd2d9;
    1230: romdata_int <= 'h72a1;
    1231: romdata_int <= 'h3b49;
    1232: romdata_int <= 'h46c; // Line Descriptor
    1233: romdata_int <= 'hab32;
    1234: romdata_int <= 'h4a6b;
    1235: romdata_int <= 'h2eb8;
    1236: romdata_int <= 'h46c; // Line Descriptor
    1237: romdata_int <= 'hb3a;
    1238: romdata_int <= 'hae48;
    1239: romdata_int <= 'h7f37;
    1240: romdata_int <= 'h46c; // Line Descriptor
    1241: romdata_int <= 'ha6b9;
    1242: romdata_int <= 'h4706;
    1243: romdata_int <= 'h1463;
    1244: romdata_int <= 'h46c; // Line Descriptor
    1245: romdata_int <= 'h267a;
    1246: romdata_int <= 'h5ec3;
    1247: romdata_int <= 'h56ca;
    1248: romdata_int <= 'h46c; // Line Descriptor
    1249: romdata_int <= 'h5828;
    1250: romdata_int <= 'h4320;
    1251: romdata_int <= 'h682c;
    1252: romdata_int <= 'h46c; // Line Descriptor
    1253: romdata_int <= 'h9a33;
    1254: romdata_int <= 'hba12;
    1255: romdata_int <= 'h9c2c;
    1256: romdata_int <= 'h56c; // Line Descriptor
    1257: romdata_int <= 'h11c;
    1258: romdata_int <= 'h9e9c;
    1259: romdata_int <= 'h889;
    1260: romdata_int <= 'he5a; // Line Descriptor
    1261: romdata_int <= 'h6c00;
    1262: romdata_int <= 'h6067;
    1263: romdata_int <= 'ha49f;
    1264: romdata_int <= 'h2b32;
    1265: romdata_int <= 'hb32a;
    1266: romdata_int <= 'h6271;
    1267: romdata_int <= 'h1c1c;
    1268: romdata_int <= 'h5e5f;
    1269: romdata_int <= 'he5a; // Line Descriptor
    1270: romdata_int <= 'h7e50;
    1271: romdata_int <= 'h6e00;
    1272: romdata_int <= 'h5a33;
    1273: romdata_int <= 'h141c;
    1274: romdata_int <= 'h6538;
    1275: romdata_int <= 'h8d08;
    1276: romdata_int <= 'h6628;
    1277: romdata_int <= 'h7e21;
    1278: romdata_int <= 'he5a; // Line Descriptor
    1279: romdata_int <= 'h7000;
    1280: romdata_int <= 'h8f12;
    1281: romdata_int <= 'h706;
    1282: romdata_int <= 'h3521;
    1283: romdata_int <= 'h26c0;
    1284: romdata_int <= 'ha03f;
    1285: romdata_int <= 'h9008;
    1286: romdata_int <= 'h9e65;
    1287: romdata_int <= 'he5a; // Line Descriptor
    1288: romdata_int <= 'h7200;
    1289: romdata_int <= 'h6640;
    1290: romdata_int <= 'h6d22;
    1291: romdata_int <= 'h2ecf;
    1292: romdata_int <= 'h3e80;
    1293: romdata_int <= 'h72ab;
    1294: romdata_int <= 'ha98;
    1295: romdata_int <= 'h80b4;
    1296: romdata_int <= 'he5a; // Line Descriptor
    1297: romdata_int <= 'h7400;
    1298: romdata_int <= 'h148c;
    1299: romdata_int <= 'he7e;
    1300: romdata_int <= 'h753f;
    1301: romdata_int <= 'h41f;
    1302: romdata_int <= 'h3023;
    1303: romdata_int <= 'h3f46;
    1304: romdata_int <= 'h4a90;
    1305: romdata_int <= 'he5a; // Line Descriptor
    1306: romdata_int <= 'h7600;
    1307: romdata_int <= 'h62ba;
    1308: romdata_int <= 'hb0b1;
    1309: romdata_int <= 'h3aee;
    1310: romdata_int <= 'h5a44;
    1311: romdata_int <= 'h68eb;
    1312: romdata_int <= 'h14b0;
    1313: romdata_int <= 'h4823;
    1314: romdata_int <= 'he5a; // Line Descriptor
    1315: romdata_int <= 'h7800;
    1316: romdata_int <= 'h7158;
    1317: romdata_int <= 'h3aee;
    1318: romdata_int <= 'h88c3;
    1319: romdata_int <= 'h645;
    1320: romdata_int <= 'h2087;
    1321: romdata_int <= 'h6c5c;
    1322: romdata_int <= 'h40ca;
    1323: romdata_int <= 'he5a; // Line Descriptor
    1324: romdata_int <= 'h7a00;
    1325: romdata_int <= 'h84fd;
    1326: romdata_int <= 'ha69d;
    1327: romdata_int <= 'h9a7d;
    1328: romdata_int <= 'h5c41;
    1329: romdata_int <= 'hb007;
    1330: romdata_int <= 'h3682;
    1331: romdata_int <= 'h4c67;
    1332: romdata_int <= 'he5a; // Line Descriptor
    1333: romdata_int <= 'h7c00;
    1334: romdata_int <= 'h2a17;
    1335: romdata_int <= 'h1715;
    1336: romdata_int <= 'had4c;
    1337: romdata_int <= 'h6d06;
    1338: romdata_int <= 'h1a64;
    1339: romdata_int <= 'h22ad;
    1340: romdata_int <= 'h583c;
    1341: romdata_int <= 'he5a; // Line Descriptor
    1342: romdata_int <= 'h7e00;
    1343: romdata_int <= 'h86f6;
    1344: romdata_int <= 'h2e2c;
    1345: romdata_int <= 'h94bb;
    1346: romdata_int <= 'h93d;
    1347: romdata_int <= 'haaed;
    1348: romdata_int <= 'h9531;
    1349: romdata_int <= 'ha51f;
    1350: romdata_int <= 'he5a; // Line Descriptor
    1351: romdata_int <= 'h8000;
    1352: romdata_int <= 'h4b1d;
    1353: romdata_int <= 'h232;
    1354: romdata_int <= 'h6af6;
    1355: romdata_int <= 'haaa2;
    1356: romdata_int <= 'h4ca4;
    1357: romdata_int <= 'h60b3;
    1358: romdata_int <= 'h23d;
    1359: romdata_int <= 'he5a; // Line Descriptor
    1360: romdata_int <= 'h8200;
    1361: romdata_int <= 'h2832;
    1362: romdata_int <= 'ha8bd;
    1363: romdata_int <= 'haf03;
    1364: romdata_int <= 'h442f;
    1365: romdata_int <= 'h64f8;
    1366: romdata_int <= 'h2abc;
    1367: romdata_int <= 'h20ef;
    1368: romdata_int <= 'he5a; // Line Descriptor
    1369: romdata_int <= 'h8400;
    1370: romdata_int <= 'h6474;
    1371: romdata_int <= 'h7c44;
    1372: romdata_int <= 'h7967;
    1373: romdata_int <= 'h726a;
    1374: romdata_int <= 'h7b56;
    1375: romdata_int <= 'h4520;
    1376: romdata_int <= 'h7c1e;
    1377: romdata_int <= 'he5a; // Line Descriptor
    1378: romdata_int <= 'h8600;
    1379: romdata_int <= 'h8cf5;
    1380: romdata_int <= 'hafe;
    1381: romdata_int <= 'ha14b;
    1382: romdata_int <= 'h36a8;
    1383: romdata_int <= 'h9c97;
    1384: romdata_int <= 'h1ea6;
    1385: romdata_int <= 'h82d5;
    1386: romdata_int <= 'he5a; // Line Descriptor
    1387: romdata_int <= 'h8800;
    1388: romdata_int <= 'h3a4a;
    1389: romdata_int <= 'h60cc;
    1390: romdata_int <= 'h98cb;
    1391: romdata_int <= 'h246e;
    1392: romdata_int <= 'hd1e;
    1393: romdata_int <= 'h563c;
    1394: romdata_int <= 'h46e5;
    1395: romdata_int <= 'he5a; // Line Descriptor
    1396: romdata_int <= 'h8a00;
    1397: romdata_int <= 'h194d;
    1398: romdata_int <= 'h268b;
    1399: romdata_int <= 'hb099;
    1400: romdata_int <= 'h8434;
    1401: romdata_int <= 'h5151;
    1402: romdata_int <= 'h426f;
    1403: romdata_int <= 'h9d13;
    1404: romdata_int <= 'he5a; // Line Descriptor
    1405: romdata_int <= 'h8c00;
    1406: romdata_int <= 'h40e;
    1407: romdata_int <= 'h5537;
    1408: romdata_int <= 'h114c;
    1409: romdata_int <= 'h1a91;
    1410: romdata_int <= 'h70b;
    1411: romdata_int <= 'ha2f3;
    1412: romdata_int <= 'h4257;
    1413: romdata_int <= 'he5a; // Line Descriptor
    1414: romdata_int <= 'h8e00;
    1415: romdata_int <= 'h3049;
    1416: romdata_int <= 'h4149;
    1417: romdata_int <= 'h535d;
    1418: romdata_int <= 'h8ea4;
    1419: romdata_int <= 'h7669;
    1420: romdata_int <= 'h8267;
    1421: romdata_int <= 'h695e;
    1422: romdata_int <= 'he5a; // Line Descriptor
    1423: romdata_int <= 'h9000;
    1424: romdata_int <= 'h100f;
    1425: romdata_int <= 'h8047;
    1426: romdata_int <= 'h92b8;
    1427: romdata_int <= 'h1ce2;
    1428: romdata_int <= 'h3911;
    1429: romdata_int <= 'ha806;
    1430: romdata_int <= 'h5a3a;
    1431: romdata_int <= 'he5a; // Line Descriptor
    1432: romdata_int <= 'h9200;
    1433: romdata_int <= 'hb2d8;
    1434: romdata_int <= 'h3203;
    1435: romdata_int <= 'h16c8;
    1436: romdata_int <= 'h2822;
    1437: romdata_int <= 'h5894;
    1438: romdata_int <= 'h2c59;
    1439: romdata_int <= 'h2eaa;
    1440: romdata_int <= 'he5a; // Line Descriptor
    1441: romdata_int <= 'h9400;
    1442: romdata_int <= 'h1685;
    1443: romdata_int <= 'h8c10;
    1444: romdata_int <= 'h5058;
    1445: romdata_int <= 'h54ee;
    1446: romdata_int <= 'h4e65;
    1447: romdata_int <= 'h3c7e;
    1448: romdata_int <= 'h31e;
    1449: romdata_int <= 'he5a; // Line Descriptor
    1450: romdata_int <= 'h9600;
    1451: romdata_int <= 'hc67;
    1452: romdata_int <= 'h5d49;
    1453: romdata_int <= 'h5632;
    1454: romdata_int <= 'h1355;
    1455: romdata_int <= 'h48e5;
    1456: romdata_int <= 'h66f3;
    1457: romdata_int <= 'h7937;
    1458: romdata_int <= 'he5a; // Line Descriptor
    1459: romdata_int <= 'h9800;
    1460: romdata_int <= 'h5ab1;
    1461: romdata_int <= 'h951c;
    1462: romdata_int <= 'h3c3d;
    1463: romdata_int <= 'h8b59;
    1464: romdata_int <= 'h4698;
    1465: romdata_int <= 'h9ef3;
    1466: romdata_int <= 'h96d9;
    1467: romdata_int <= 'he5a; // Line Descriptor
    1468: romdata_int <= 'h9a00;
    1469: romdata_int <= 'h74cf;
    1470: romdata_int <= 'h2433;
    1471: romdata_int <= 'h9760;
    1472: romdata_int <= 'h1f4f;
    1473: romdata_int <= 'h6a91;
    1474: romdata_int <= 'hac76;
    1475: romdata_int <= 'h8144;
    1476: romdata_int <= 'he5a; // Line Descriptor
    1477: romdata_int <= 'h9c00;
    1478: romdata_int <= 'h8ef;
    1479: romdata_int <= 'h9b00;
    1480: romdata_int <= 'ha88;
    1481: romdata_int <= 'h3321;
    1482: romdata_int <= 'h855f;
    1483: romdata_int <= 'h8f1c;
    1484: romdata_int <= 'h1355;
    1485: romdata_int <= 'he5a; // Line Descriptor
    1486: romdata_int <= 'h9e00;
    1487: romdata_int <= 'h586b;
    1488: romdata_int <= 'h4915;
    1489: romdata_int <= 'h6f5b;
    1490: romdata_int <= 'h394c;
    1491: romdata_int <= 'h40bd;
    1492: romdata_int <= 'h2511;
    1493: romdata_int <= 'haf61;
    1494: romdata_int <= 'he5a; // Line Descriptor
    1495: romdata_int <= 'ha000;
    1496: romdata_int <= 'h98f2;
    1497: romdata_int <= 'h7334;
    1498: romdata_int <= 'h4f4c;
    1499: romdata_int <= 'h12c;
    1500: romdata_int <= 'h5ea5;
    1501: romdata_int <= 'h8a7e;
    1502: romdata_int <= 'h184f;
    1503: romdata_int <= 'he5a; // Line Descriptor
    1504: romdata_int <= 'ha200;
    1505: romdata_int <= 'h934a;
    1506: romdata_int <= 'h103;
    1507: romdata_int <= 'ha602;
    1508: romdata_int <= 'h2236;
    1509: romdata_int <= 'h53e;
    1510: romdata_int <= 'h32e4;
    1511: romdata_int <= 'h54f5;
    1512: romdata_int <= 'he5a; // Line Descriptor
    1513: romdata_int <= 'ha400;
    1514: romdata_int <= 'h46ad;
    1515: romdata_int <= 'h8e3e;
    1516: romdata_int <= 'ha8f2;
    1517: romdata_int <= 'he2c;
    1518: romdata_int <= 'h26a0;
    1519: romdata_int <= 'h9afc;
    1520: romdata_int <= 'h70b0;
    1521: romdata_int <= 'he5a; // Line Descriptor
    1522: romdata_int <= 'ha600;
    1523: romdata_int <= 'hab4e;
    1524: romdata_int <= 'h6213;
    1525: romdata_int <= 'h7670;
    1526: romdata_int <= 'h7f44;
    1527: romdata_int <= 'h9921;
    1528: romdata_int <= 'h3475;
    1529: romdata_int <= 'h7438;
    1530: romdata_int <= 'he5a; // Line Descriptor
    1531: romdata_int <= 'ha800;
    1532: romdata_int <= 'had1;
    1533: romdata_int <= 'h1eb8;
    1534: romdata_int <= 'h7020;
    1535: romdata_int <= 'h870f;
    1536: romdata_int <= 'h1129;
    1537: romdata_int <= 'h43;
    1538: romdata_int <= 'h6e05;
    1539: romdata_int <= 'he5a; // Line Descriptor
    1540: romdata_int <= 'haa00;
    1541: romdata_int <= 'had50;
    1542: romdata_int <= 'h88f7;
    1543: romdata_int <= 'h2d32;
    1544: romdata_int <= 'h7adf;
    1545: romdata_int <= 'h2925;
    1546: romdata_int <= 'h4a45;
    1547: romdata_int <= 'h5313;
    1548: romdata_int <= 'he5a; // Line Descriptor
    1549: romdata_int <= 'hac00;
    1550: romdata_int <= 'h380a;
    1551: romdata_int <= 'had44;
    1552: romdata_int <= 'hcec;
    1553: romdata_int <= 'h8c89;
    1554: romdata_int <= 'h16aa;
    1555: romdata_int <= 'hb366;
    1556: romdata_int <= 'h88ce;
    1557: romdata_int <= 'he5a; // Line Descriptor
    1558: romdata_int <= 'hae00;
    1559: romdata_int <= 'h80e1;
    1560: romdata_int <= 'haa42;
    1561: romdata_int <= 'h6328;
    1562: romdata_int <= 'h18b5;
    1563: romdata_int <= 'h5c19;
    1564: romdata_int <= 'h824;
    1565: romdata_int <= 'ha6d9;
    1566: romdata_int <= 'he5a; // Line Descriptor
    1567: romdata_int <= 'hb000;
    1568: romdata_int <= 'h3645;
    1569: romdata_int <= 'h7e84;
    1570: romdata_int <= 'ha2fd;
    1571: romdata_int <= 'h90ad;
    1572: romdata_int <= 'hf09;
    1573: romdata_int <= 'ha4a7;
    1574: romdata_int <= 'h86e8;
    1575: romdata_int <= 'he5a; // Line Descriptor
    1576: romdata_int <= 'hb200;
    1577: romdata_int <= 'h4325;
    1578: romdata_int <= 'h7517;
    1579: romdata_int <= 'h60d3;
    1580: romdata_int <= 'h30cc;
    1581: romdata_int <= 'h7c62;
    1582: romdata_int <= 'h3a8d;
    1583: romdata_int <= 'h924e;
    1584: romdata_int <= 'h45a; // Line Descriptor
    1585: romdata_int <= 'h0;
    1586: romdata_int <= 'h9aa1;
    1587: romdata_int <= 'h4715;
    1588: romdata_int <= 'h45a; // Line Descriptor
    1589: romdata_int <= 'h200;
    1590: romdata_int <= 'h4c2b;
    1591: romdata_int <= 'h1401;
    1592: romdata_int <= 'h45a; // Line Descriptor
    1593: romdata_int <= 'h400;
    1594: romdata_int <= 'h2672;
    1595: romdata_int <= 'h7802;
    1596: romdata_int <= 'h45a; // Line Descriptor
    1597: romdata_int <= 'h600;
    1598: romdata_int <= 'h910b;
    1599: romdata_int <= 'h5808;
    1600: romdata_int <= 'h45a; // Line Descriptor
    1601: romdata_int <= 'h800;
    1602: romdata_int <= 'h6a89;
    1603: romdata_int <= 'h422e;
    1604: romdata_int <= 'h45a; // Line Descriptor
    1605: romdata_int <= 'ha00;
    1606: romdata_int <= 'h29a;
    1607: romdata_int <= 'h9cb0;
    1608: romdata_int <= 'h45a; // Line Descriptor
    1609: romdata_int <= 'hc00;
    1610: romdata_int <= 'haeec;
    1611: romdata_int <= 'h700b;
    1612: romdata_int <= 'h45a; // Line Descriptor
    1613: romdata_int <= 'he00;
    1614: romdata_int <= 'h883a;
    1615: romdata_int <= 'hb2a1;
    1616: romdata_int <= 'h45a; // Line Descriptor
    1617: romdata_int <= 'h1000;
    1618: romdata_int <= 'h9d38;
    1619: romdata_int <= 'h7659;
    1620: romdata_int <= 'h45a; // Line Descriptor
    1621: romdata_int <= 'h1200;
    1622: romdata_int <= 'h2eb8;
    1623: romdata_int <= 'h387b;
    1624: romdata_int <= 'h45a; // Line Descriptor
    1625: romdata_int <= 'h1400;
    1626: romdata_int <= 'h3eb9;
    1627: romdata_int <= 'h1b3b;
    1628: romdata_int <= 'h45a; // Line Descriptor
    1629: romdata_int <= 'h1600;
    1630: romdata_int <= 'h3c9b;
    1631: romdata_int <= 'h8312;
    1632: romdata_int <= 'h45a; // Line Descriptor
    1633: romdata_int <= 'h1800;
    1634: romdata_int <= 'h4f65;
    1635: romdata_int <= 'h9ec7;
    1636: romdata_int <= 'h45a; // Line Descriptor
    1637: romdata_int <= 'h1a00;
    1638: romdata_int <= 'h2279;
    1639: romdata_int <= 'h861e;
    1640: romdata_int <= 'h45a; // Line Descriptor
    1641: romdata_int <= 'h1c00;
    1642: romdata_int <= 'h5eef;
    1643: romdata_int <= 'h4c2a;
    1644: romdata_int <= 'h45a; // Line Descriptor
    1645: romdata_int <= 'h1e00;
    1646: romdata_int <= 'h4928;
    1647: romdata_int <= 'h48a;
    1648: romdata_int <= 'h45a; // Line Descriptor
    1649: romdata_int <= 'h2000;
    1650: romdata_int <= 'h3455;
    1651: romdata_int <= 'h3061;
    1652: romdata_int <= 'h45a; // Line Descriptor
    1653: romdata_int <= 'h2200;
    1654: romdata_int <= 'h6ea5;
    1655: romdata_int <= 'h90e0;
    1656: romdata_int <= 'h45a; // Line Descriptor
    1657: romdata_int <= 'h2400;
    1658: romdata_int <= 'h76ae;
    1659: romdata_int <= 'h9911;
    1660: romdata_int <= 'h45a; // Line Descriptor
    1661: romdata_int <= 'h2600;
    1662: romdata_int <= 'ha562;
    1663: romdata_int <= 'h4e5f;
    1664: romdata_int <= 'h45a; // Line Descriptor
    1665: romdata_int <= 'h2800;
    1666: romdata_int <= 'hb0dd;
    1667: romdata_int <= 'h232e;
    1668: romdata_int <= 'h45a; // Line Descriptor
    1669: romdata_int <= 'h2a00;
    1670: romdata_int <= 'h792c;
    1671: romdata_int <= 'h52a7;
    1672: romdata_int <= 'h45a; // Line Descriptor
    1673: romdata_int <= 'h2c00;
    1674: romdata_int <= 'h5243;
    1675: romdata_int <= 'h1328;
    1676: romdata_int <= 'h45a; // Line Descriptor
    1677: romdata_int <= 'h2e00;
    1678: romdata_int <= 'h5673;
    1679: romdata_int <= 'h207c;
    1680: romdata_int <= 'h45a; // Line Descriptor
    1681: romdata_int <= 'h3000;
    1682: romdata_int <= 'h726a;
    1683: romdata_int <= 'h6494;
    1684: romdata_int <= 'h45a; // Line Descriptor
    1685: romdata_int <= 'h3200;
    1686: romdata_int <= 'h7a4e;
    1687: romdata_int <= 'h4ac4;
    1688: romdata_int <= 'h45a; // Line Descriptor
    1689: romdata_int <= 'h3400;
    1690: romdata_int <= 'ha60f;
    1691: romdata_int <= 'h92d8;
    1692: romdata_int <= 'h45a; // Line Descriptor
    1693: romdata_int <= 'h3600;
    1694: romdata_int <= 'h1f2b;
    1695: romdata_int <= 'h1c64;
    1696: romdata_int <= 'h45a; // Line Descriptor
    1697: romdata_int <= 'h3800;
    1698: romdata_int <= 'h40d5;
    1699: romdata_int <= 'ha062;
    1700: romdata_int <= 'h45a; // Line Descriptor
    1701: romdata_int <= 'h3a00;
    1702: romdata_int <= 'h7cc9;
    1703: romdata_int <= 'h5f54;
    1704: romdata_int <= 'h45a; // Line Descriptor
    1705: romdata_int <= 'h3c00;
    1706: romdata_int <= 'h1ae7;
    1707: romdata_int <= 'h3613;
    1708: romdata_int <= 'h45a; // Line Descriptor
    1709: romdata_int <= 'h3e00;
    1710: romdata_int <= 'h1c83;
    1711: romdata_int <= 'h2b18;
    1712: romdata_int <= 'h45a; // Line Descriptor
    1713: romdata_int <= 'h4000;
    1714: romdata_int <= 'h760;
    1715: romdata_int <= 'h6ac5;
    1716: romdata_int <= 'h45a; // Line Descriptor
    1717: romdata_int <= 'h4200;
    1718: romdata_int <= 'ha949;
    1719: romdata_int <= 'h9667;
    1720: romdata_int <= 'h45a; // Line Descriptor
    1721: romdata_int <= 'h4400;
    1722: romdata_int <= 'h5088;
    1723: romdata_int <= 'h7b27;
    1724: romdata_int <= 'h45a; // Line Descriptor
    1725: romdata_int <= 'h4600;
    1726: romdata_int <= 'h5c48;
    1727: romdata_int <= 'h2d22;
    1728: romdata_int <= 'h45a; // Line Descriptor
    1729: romdata_int <= 'h4800;
    1730: romdata_int <= 'h8322;
    1731: romdata_int <= 'ha27c;
    1732: romdata_int <= 'h45a; // Line Descriptor
    1733: romdata_int <= 'h4a00;
    1734: romdata_int <= 'h2055;
    1735: romdata_int <= 'h692b;
    1736: romdata_int <= 'h45a; // Line Descriptor
    1737: romdata_int <= 'h4c00;
    1738: romdata_int <= 'hb5;
    1739: romdata_int <= 'h285e;
    1740: romdata_int <= 'h45a; // Line Descriptor
    1741: romdata_int <= 'h4e00;
    1742: romdata_int <= 'h9482;
    1743: romdata_int <= 'h5070;
    1744: romdata_int <= 'h45a; // Line Descriptor
    1745: romdata_int <= 'h5000;
    1746: romdata_int <= 'ha34d;
    1747: romdata_int <= 'hd52;
    1748: romdata_int <= 'h45a; // Line Descriptor
    1749: romdata_int <= 'h5200;
    1750: romdata_int <= 'h960e;
    1751: romdata_int <= 'h44ab;
    1752: romdata_int <= 'h45a; // Line Descriptor
    1753: romdata_int <= 'h5400;
    1754: romdata_int <= 'h324c;
    1755: romdata_int <= 'h18c5;
    1756: romdata_int <= 'h45a; // Line Descriptor
    1757: romdata_int <= 'h5600;
    1758: romdata_int <= 'h1361;
    1759: romdata_int <= 'h8a8a;
    1760: romdata_int <= 'h45a; // Line Descriptor
    1761: romdata_int <= 'h5800;
    1762: romdata_int <= 'ha164;
    1763: romdata_int <= 'h3ee9;
    1764: romdata_int <= 'h45a; // Line Descriptor
    1765: romdata_int <= 'h5a00;
    1766: romdata_int <= 'h24a1;
    1767: romdata_int <= 'h844d;
    1768: romdata_int <= 'h45a; // Line Descriptor
    1769: romdata_int <= 'h5c00;
    1770: romdata_int <= 'h9e0a;
    1771: romdata_int <= 'h916;
    1772: romdata_int <= 'h45a; // Line Descriptor
    1773: romdata_int <= 'h5e00;
    1774: romdata_int <= 'h6c32;
    1775: romdata_int <= 'h34f3;
    1776: romdata_int <= 'h45a; // Line Descriptor
    1777: romdata_int <= 'h6000;
    1778: romdata_int <= 'h8a58;
    1779: romdata_int <= 'haef1;
    1780: romdata_int <= 'h45a; // Line Descriptor
    1781: romdata_int <= 'h6200;
    1782: romdata_int <= 'h2c37;
    1783: romdata_int <= 'h66e5;
    1784: romdata_int <= 'h45a; // Line Descriptor
    1785: romdata_int <= 'h6400;
    1786: romdata_int <= 'h5449;
    1787: romdata_int <= 'h3c1e;
    1788: romdata_int <= 'h45a; // Line Descriptor
    1789: romdata_int <= 'h6600;
    1790: romdata_int <= 'h688d;
    1791: romdata_int <= 'h1031;
    1792: romdata_int <= 'h45a; // Line Descriptor
    1793: romdata_int <= 'h6800;
    1794: romdata_int <= 'h4544;
    1795: romdata_int <= 'h6e06;
    1796: romdata_int <= 'h55a; // Line Descriptor
    1797: romdata_int <= 'h6a00;
    1798: romdata_int <= 'hed6;
    1799: romdata_int <= 'h56df;
    1800: romdata_int <= 'h1648; // Line Descriptor
    1801: romdata_int <= 'h3d37;
    1802: romdata_int <= 'h748e;
    1803: romdata_int <= 'h44a1;
    1804: romdata_int <= 'h6b15;
    1805: romdata_int <= 'h29b;
    1806: romdata_int <= 'h5428;
    1807: romdata_int <= 'h342b;
    1808: romdata_int <= 'h3601;
    1809: romdata_int <= 'h124e;
    1810: romdata_int <= 'hed;
    1811: romdata_int <= 'h7c72;
    1812: romdata_int <= 'h4602;
    1813: romdata_int <= 'h1648; // Line Descriptor
    1814: romdata_int <= 'h3f5c;
    1815: romdata_int <= 'h24e1;
    1816: romdata_int <= 'h2eec;
    1817: romdata_int <= 'h480b;
    1818: romdata_int <= 'h3316;
    1819: romdata_int <= 'h3164;
    1820: romdata_int <= 'h143a;
    1821: romdata_int <= 'h4aa1;
    1822: romdata_int <= 'h7f39;
    1823: romdata_int <= 'h32f0;
    1824: romdata_int <= 'h6738;
    1825: romdata_int <= 'h6e59;
    1826: romdata_int <= 'h1648; // Line Descriptor
    1827: romdata_int <= 'h4299;
    1828: romdata_int <= 'h3b3d;
    1829: romdata_int <= 'h565;
    1830: romdata_int <= 'h78c7;
    1831: romdata_int <= 'h384c;
    1832: romdata_int <= 'h2b0b;
    1833: romdata_int <= 'h2879;
    1834: romdata_int <= 'h221e;
    1835: romdata_int <= 'h26bc;
    1836: romdata_int <= 'h549d;
    1837: romdata_int <= 'h72ef;
    1838: romdata_int <= 'h5a2a;
    1839: romdata_int <= 'h1648; // Line Descriptor
    1840: romdata_int <= 'h2ae6;
    1841: romdata_int <= 'h6334;
    1842: romdata_int <= 'h46ae;
    1843: romdata_int <= 'h7b11;
    1844: romdata_int <= 'h4347;
    1845: romdata_int <= 'h46a0;
    1846: romdata_int <= 'h1162;
    1847: romdata_int <= 'h1a5f;
    1848: romdata_int <= 'h7760;
    1849: romdata_int <= 'h4448;
    1850: romdata_int <= 'h1add;
    1851: romdata_int <= 'h2d2e;
    1852: romdata_int <= 'h1648; // Line Descriptor
    1853: romdata_int <= 'h52e5;
    1854: romdata_int <= 'h1ec9;
    1855: romdata_int <= 'h166a;
    1856: romdata_int <= 'h7694;
    1857: romdata_int <= 'h24f2;
    1858: romdata_int <= 'h3e9a;
    1859: romdata_int <= 'h7e4e;
    1860: romdata_int <= 'h56c4;
    1861: romdata_int <= 'h2b50;
    1862: romdata_int <= 'h6123;
    1863: romdata_int <= 'h480f;
    1864: romdata_int <= 'h88d8;
    1865: romdata_int <= 'h1648; // Line Descriptor
    1866: romdata_int <= 'h184a;
    1867: romdata_int <= 'h8877;
    1868: romdata_int <= 'h7ae7;
    1869: romdata_int <= 'h8413;
    1870: romdata_int <= 'h264e;
    1871: romdata_int <= 'h485a;
    1872: romdata_int <= 'h6483;
    1873: romdata_int <= 'h3b18;
    1874: romdata_int <= 'h740e;
    1875: romdata_int <= 'h4ad0;
    1876: romdata_int <= 'h2360;
    1877: romdata_int <= 'h76c5;
    1878: romdata_int <= 'h1648; // Line Descriptor
    1879: romdata_int <= 'h501;
    1880: romdata_int <= 'h7934;
    1881: romdata_int <= 'h4122;
    1882: romdata_int <= 'h307c;
    1883: romdata_int <= 'h2a4b;
    1884: romdata_int <= 'h86d9;
    1885: romdata_int <= 'hc55;
    1886: romdata_int <= 'h872b;
    1887: romdata_int <= 'h8806;
    1888: romdata_int <= 'h805f;
    1889: romdata_int <= 'h36b5;
    1890: romdata_int <= 'h445e;
    1891: romdata_int <= 'h1648; // Line Descriptor
    1892: romdata_int <= 'h1275;
    1893: romdata_int <= 'h1c41;
    1894: romdata_int <= 'h684c;
    1895: romdata_int <= 'h40c5;
    1896: romdata_int <= 'h1a33;
    1897: romdata_int <= 'h8311;
    1898: romdata_int <= 'h961;
    1899: romdata_int <= 'h28a;
    1900: romdata_int <= 'h6b4a;
    1901: romdata_int <= 'h5e7d;
    1902: romdata_int <= 'h2764;
    1903: romdata_int <= 'h64e9;
    1904: romdata_int <= 'h1648; // Line Descriptor
    1905: romdata_int <= 'h592a;
    1906: romdata_int <= 'h5d58;
    1907: romdata_int <= 'h1058;
    1908: romdata_int <= 'h3cf1;
    1909: romdata_int <= 'h1062;
    1910: romdata_int <= 'h42c1;
    1911: romdata_int <= 'h5837;
    1912: romdata_int <= 'h80e5;
    1913: romdata_int <= 'h4b2;
    1914: romdata_int <= 'h1079;
    1915: romdata_int <= 'h3c49;
    1916: romdata_int <= 'h5c1e;
    1917: romdata_int <= 'h1648; // Line Descriptor
    1918: romdata_int <= 'h6b38;
    1919: romdata_int <= 'h6a21;
    1920: romdata_int <= 'h7308;
    1921: romdata_int <= 'h5228;
    1922: romdata_int <= 'h172c;
    1923: romdata_int <= 'h21a;
    1924: romdata_int <= 'h2668;
    1925: romdata_int <= 'h5a4e;
    1926: romdata_int <= 'h4d3f;
    1927: romdata_int <= 'h2141;
    1928: romdata_int <= 'h2f1d;
    1929: romdata_int <= 'h6312;
    1930: romdata_int <= 'h1648; // Line Descriptor
    1931: romdata_int <= 'h5418;
    1932: romdata_int <= 'h3840;
    1933: romdata_int <= 'h2922;
    1934: romdata_int <= 'h36cf;
    1935: romdata_int <= 'h3e80;
    1936: romdata_int <= 'h38ab;
    1937: romdata_int <= 'h8098;
    1938: romdata_int <= 'hcb4;
    1939: romdata_int <= 'he3e;
    1940: romdata_int <= 'h8625;
    1941: romdata_int <= 'h3ae4;
    1942: romdata_int <= 'h8e0a;
    1943: romdata_int <= 'h1648; // Line Descriptor
    1944: romdata_int <= 'h165c;
    1945: romdata_int <= 'h18ca;
    1946: romdata_int <= 'h306;
    1947: romdata_int <= 'h3b37;
    1948: romdata_int <= 'h2933;
    1949: romdata_int <= 'h32b0;
    1950: romdata_int <= 'h1688;
    1951: romdata_int <= 'h8b61;
    1952: romdata_int <= 'h506b;
    1953: romdata_int <= 'h4cfd;
    1954: romdata_int <= 'h129d;
    1955: romdata_int <= 'h87d;
    1956: romdata_int <= 'h1648; // Line Descriptor
    1957: romdata_int <= 'h4d15;
    1958: romdata_int <= 'h774c;
    1959: romdata_int <= 'h6106;
    1960: romdata_int <= 'hc64;
    1961: romdata_int <= 'h58ad;
    1962: romdata_int <= 'h7c3c;
    1963: romdata_int <= 'h6716;
    1964: romdata_int <= 'h7255;
    1965: romdata_int <= 'h6f23;
    1966: romdata_int <= 'h5610;
    1967: romdata_int <= 'h747;
    1968: romdata_int <= 'h8b58;
    1969: romdata_int <= 'h1648; // Line Descriptor
    1970: romdata_int <= 'h480a;
    1971: romdata_int <= 'h8c9a;
    1972: romdata_int <= 'h3ccb;
    1973: romdata_int <= 'h1d1d;
    1974: romdata_int <= 'h5e32;
    1975: romdata_int <= 'h20f6;
    1976: romdata_int <= 'h18a2;
    1977: romdata_int <= 'h46a4;
    1978: romdata_int <= 'h62b3;
    1979: romdata_int <= 'h143d;
    1980: romdata_int <= 'h6a72;
    1981: romdata_int <= 'h613e;
    1982: romdata_int <= 'h1648; // Line Descriptor
    1983: romdata_int <= 'h2481;
    1984: romdata_int <= 'h434d;
    1985: romdata_int <= 'h88b;
    1986: romdata_int <= 'h8299;
    1987: romdata_int <= 'h434;
    1988: romdata_int <= 'h7b51;
    1989: romdata_int <= 'h886f;
    1990: romdata_int <= 'h3513;
    1991: romdata_int <= 'h640b;
    1992: romdata_int <= 'h687a;
    1993: romdata_int <= 'h2428;
    1994: romdata_int <= 'h6645;
    1995: romdata_int <= 'h1648; // Line Descriptor
    1996: romdata_int <= 'h1e69;
    1997: romdata_int <= 'h4e67;
    1998: romdata_int <= 'h595e;
    1999: romdata_int <= 'h7041;
    2000: romdata_int <= 'hc8;
    2001: romdata_int <= 'h1b3f;
    2002: romdata_int <= 'h8e4c;
    2003: romdata_int <= 'h1c6f;
    2004: romdata_int <= 'h1750;
    2005: romdata_int <= 'h2ab5;
    2006: romdata_int <= 'h500f;
    2007: romdata_int <= 'h2047;
    2008: romdata_int <= 'h1648; // Line Descriptor
    2009: romdata_int <= 'h3430;
    2010: romdata_int <= 'h6c80;
    2011: romdata_int <= 'h36b5;
    2012: romdata_int <= 'h72db;
    2013: romdata_int <= 'h4a67;
    2014: romdata_int <= 'h7749;
    2015: romdata_int <= 'h7032;
    2016: romdata_int <= 'h4355;
    2017: romdata_int <= 'h6ce5;
    2018: romdata_int <= 'h16f3;
    2019: romdata_int <= 'h8d37;
    2020: romdata_int <= 'h6ccb;
    2021: romdata_int <= 'h1648; // Line Descriptor
    2022: romdata_int <= 'h6d9;
    2023: romdata_int <= 'h34d4;
    2024: romdata_int <= 'h2c3a;
    2025: romdata_int <= 'h893b;
    2026: romdata_int <= 'h1451;
    2027: romdata_int <= 'h6ba;
    2028: romdata_int <= 'h1d4c;
    2029: romdata_int <= 'h82eb;
    2030: romdata_int <= 'h32cf;
    2031: romdata_int <= 'h6c33;
    2032: romdata_int <= 'hd60;
    2033: romdata_int <= 'h4b4f;
    2034: romdata_int <= 'h1648; // Line Descriptor
    2035: romdata_int <= 'h7159;
    2036: romdata_int <= 'h2ae3;
    2037: romdata_int <= 'hee4;
    2038: romdata_int <= 'h8aba;
    2039: romdata_int <= 'h6ee6;
    2040: romdata_int <= 'h5670;
    2041: romdata_int <= 'h5b57;
    2042: romdata_int <= 'h832;
    2043: romdata_int <= 'h7167;
    2044: romdata_int <= 'h879;
    2045: romdata_int <= 'h3885;
    2046: romdata_int <= 'h7b1a;
    2047: romdata_int <= 'h1648; // Line Descriptor
    2048: romdata_int <= 'h7233;
    2049: romdata_int <= 'h4aef;
    2050: romdata_int <= 'h2100;
    2051: romdata_int <= 'h8c88;
    2052: romdata_int <= 'h2f21;
    2053: romdata_int <= 'h6d5f;
    2054: romdata_int <= 'h8b1c;
    2055: romdata_int <= 'h8555;
    2056: romdata_int <= 'h44b8;
    2057: romdata_int <= 'h7646;
    2058: romdata_int <= 'h8ec4;
    2059: romdata_int <= 'h287a;
    2060: romdata_int <= 'h1648; // Line Descriptor
    2061: romdata_int <= 'h4ee4;
    2062: romdata_int <= 'hcf5;
    2063: romdata_int <= 'h50d5;
    2064: romdata_int <= 'h64fc;
    2065: romdata_int <= 'h5162;
    2066: romdata_int <= 'h6218;
    2067: romdata_int <= 'h2454;
    2068: romdata_int <= 'h4f2f;
    2069: romdata_int <= 'h58c7;
    2070: romdata_int <= 'h7aad;
    2071: romdata_int <= 'h303e;
    2072: romdata_int <= 'h84f2;
    2073: romdata_int <= 'h1648; // Line Descriptor
    2074: romdata_int <= 'h4013;
    2075: romdata_int <= 'h8e70;
    2076: romdata_int <= 'h5f44;
    2077: romdata_int <= 'h8f21;
    2078: romdata_int <= 'h6875;
    2079: romdata_int <= 'h6838;
    2080: romdata_int <= 'h60b3;
    2081: romdata_int <= 'h6162;
    2082: romdata_int <= 'h7b35;
    2083: romdata_int <= 'h2ce6;
    2084: romdata_int <= 'h8458;
    2085: romdata_int <= 'h3152;
    2086: romdata_int <= 'h1648; // Line Descriptor
    2087: romdata_int <= 'h7f5c;
    2088: romdata_int <= 'h5547;
    2089: romdata_int <= 'h7001;
    2090: romdata_int <= 'h1242;
    2091: romdata_int <= 'h691;
    2092: romdata_int <= 'h139;
    2093: romdata_int <= 'h4e77;
    2094: romdata_int <= 'h4087;
    2095: romdata_int <= 'h3d61;
    2096: romdata_int <= 'had1;
    2097: romdata_int <= 'h7019;
    2098: romdata_int <= 'h1038;
    2099: romdata_int <= 'h1648; // Line Descriptor
    2100: romdata_int <= 'h2205;
    2101: romdata_int <= 'h8125;
    2102: romdata_int <= 'h14bb;
    2103: romdata_int <= 'h664b;
    2104: romdata_int <= 'h44ee;
    2105: romdata_int <= 'h4452;
    2106: romdata_int <= 'h408e;
    2107: romdata_int <= 'h28a6;
    2108: romdata_int <= 'h2550;
    2109: romdata_int <= 'h62f7;
    2110: romdata_int <= 'h1f32;
    2111: romdata_int <= 'h68df;
    2112: romdata_int <= 'h1648; // Line Descriptor
    2113: romdata_int <= 'h56b5;
    2114: romdata_int <= 'h86;
    2115: romdata_int <= 'h8554;
    2116: romdata_int <= 'h5cb6;
    2117: romdata_int <= 'h474b;
    2118: romdata_int <= 'h4a65;
    2119: romdata_int <= 'h8d12;
    2120: romdata_int <= 'h4829;
    2121: romdata_int <= 'h14ea;
    2122: romdata_int <= 'h243;
    2123: romdata_int <= 'h5d4c;
    2124: romdata_int <= 'had2;
    2125: romdata_int <= 'h1648; // Line Descriptor
    2126: romdata_int <= 'hd1d;
    2127: romdata_int <= 'h3231;
    2128: romdata_int <= 'haa0;
    2129: romdata_int <= 'h4d44;
    2130: romdata_int <= 'h822;
    2131: romdata_int <= 'h74f4;
    2132: romdata_int <= 'h530b;
    2133: romdata_int <= 'h1918;
    2134: romdata_int <= 'h78fa;
    2135: romdata_int <= 'h5355;
    2136: romdata_int <= 'heb8;
    2137: romdata_int <= 'h5015;
    2138: romdata_int <= 'h1648; // Line Descriptor
    2139: romdata_int <= 'h5f05;
    2140: romdata_int <= 'h4925;
    2141: romdata_int <= 'h3f17;
    2142: romdata_int <= 'h2cd3;
    2143: romdata_int <= 'h22cc;
    2144: romdata_int <= 'h5062;
    2145: romdata_int <= 'h2c8d;
    2146: romdata_int <= 'h5e4e;
    2147: romdata_int <= 'h703;
    2148: romdata_int <= 'h5911;
    2149: romdata_int <= 'h88ad;
    2150: romdata_int <= 'h82c2;
    2151: romdata_int <= 'h1648; // Line Descriptor
    2152: romdata_int <= 'h2e39;
    2153: romdata_int <= 'h2629;
    2154: romdata_int <= 'h6f3;
    2155: romdata_int <= 'h1ee2;
    2156: romdata_int <= 'h6136;
    2157: romdata_int <= 'hf2a;
    2158: romdata_int <= 'h2e6e;
    2159: romdata_int <= 'h2106;
    2160: romdata_int <= 'h2e4d;
    2161: romdata_int <= 'h6e6f;
    2162: romdata_int <= 'h4744;
    2163: romdata_int <= 'h3a5e;
    2164: romdata_int <= 'h1648; // Line Descriptor
    2165: romdata_int <= 'h8693;
    2166: romdata_int <= 'h7f53;
    2167: romdata_int <= 'h8ac6;
    2168: romdata_int <= 'h6238;
    2169: romdata_int <= 'h7464;
    2170: romdata_int <= 'h6a44;
    2171: romdata_int <= 'h7861;
    2172: romdata_int <= 'h8c0e;
    2173: romdata_int <= 'ha0b;
    2174: romdata_int <= 'h1d3e;
    2175: romdata_int <= 'h351c;
    2176: romdata_int <= 'h8c3b;
    2177: romdata_int <= 'h1648; // Line Descriptor
    2178: romdata_int <= 'h7d28;
    2179: romdata_int <= 'h6eb7;
    2180: romdata_int <= 'h233f;
    2181: romdata_int <= 'h2046;
    2182: romdata_int <= 'ha35;
    2183: romdata_int <= 'h3d49;
    2184: romdata_int <= 'h84c4;
    2185: romdata_int <= 'h548a;
    2186: romdata_int <= 'h2d08;
    2187: romdata_int <= 'h6547;
    2188: romdata_int <= 'h4e7b;
    2189: romdata_int <= 'h1d60;
    2190: romdata_int <= 'h1648; // Line Descriptor
    2191: romdata_int <= 'he56;
    2192: romdata_int <= 'h3132;
    2193: romdata_int <= 'h5a6b;
    2194: romdata_int <= 'h7cb8;
    2195: romdata_int <= 'h4e37;
    2196: romdata_int <= 'h1349;
    2197: romdata_int <= 'h3ae4;
    2198: romdata_int <= 'h393a;
    2199: romdata_int <= 'h5248;
    2200: romdata_int <= 'h5b37;
    2201: romdata_int <= 'h434f;
    2202: romdata_int <= 'h1483;
    2203: romdata_int <= 'h1648; // Line Descriptor
    2204: romdata_int <= 'h746e;
    2205: romdata_int <= 'h12a9;
    2206: romdata_int <= 'h1a28;
    2207: romdata_int <= 'h5520;
    2208: romdata_int <= 'he2c;
    2209: romdata_int <= 'ha78;
    2210: romdata_int <= 'h6ea4;
    2211: romdata_int <= 'h8f55;
    2212: romdata_int <= 'h1e8f;
    2213: romdata_int <= 'h7f65;
    2214: romdata_int <= 'h82ec;
    2215: romdata_int <= 'h2633;
    2216: romdata_int <= 'h1648; // Line Descriptor
    2217: romdata_int <= 'h331c;
    2218: romdata_int <= 'h7c9c;
    2219: romdata_int <= 'h6489;
    2220: romdata_int <= 'h7f3c;
    2221: romdata_int <= 'h6c23;
    2222: romdata_int <= 'h1e75;
    2223: romdata_int <= 'h3633;
    2224: romdata_int <= 'h3e4b;
    2225: romdata_int <= 'h159;
    2226: romdata_int <= 'h2930;
    2227: romdata_int <= 'h40df;
    2228: romdata_int <= 'h38fd;
    2229: romdata_int <= 'h1648; // Line Descriptor
    2230: romdata_int <= 'h72;
    2231: romdata_int <= 'h864f;
    2232: romdata_int <= 'h6708;
    2233: romdata_int <= 'h5a76;
    2234: romdata_int <= 'h195a;
    2235: romdata_int <= 'h5c59;
    2236: romdata_int <= 'h49c;
    2237: romdata_int <= 'h6891;
    2238: romdata_int <= 'h7ce3;
    2239: romdata_int <= 'h3e96;
    2240: romdata_int <= 'h789e;
    2241: romdata_int <= 'h286;
    2242: romdata_int <= 'h1648; // Line Descriptor
    2243: romdata_int <= 'h80e1;
    2244: romdata_int <= 'h569c;
    2245: romdata_int <= 'h535a;
    2246: romdata_int <= 'h5620;
    2247: romdata_int <= 'h86af;
    2248: romdata_int <= 'h4d0a;
    2249: romdata_int <= 'h7264;
    2250: romdata_int <= 'h5c63;
    2251: romdata_int <= 'h6758;
    2252: romdata_int <= 'h7428;
    2253: romdata_int <= 'h423;
    2254: romdata_int <= 'h1aa3;
    2255: romdata_int <= 'h1648; // Line Descriptor
    2256: romdata_int <= 'h3632;
    2257: romdata_int <= 'h8252;
    2258: romdata_int <= 'h4cc0;
    2259: romdata_int <= 'h3415;
    2260: romdata_int <= 'h8141;
    2261: romdata_int <= 'h2258;
    2262: romdata_int <= 'h5e27;
    2263: romdata_int <= 'h10f6;
    2264: romdata_int <= 'h3022;
    2265: romdata_int <= 'h1867;
    2266: romdata_int <= 'h8a07;
    2267: romdata_int <= 'h78d0;
    2268: romdata_int <= 'h448; // Line Descriptor
    2269: romdata_int <= 'h0;
    2270: romdata_int <= 'h4701;
    2271: romdata_int <= 'h1b03;
    2272: romdata_int <= 'h448; // Line Descriptor
    2273: romdata_int <= 'h200;
    2274: romdata_int <= 'h7c91;
    2275: romdata_int <= 'h6429;
    2276: romdata_int <= 'h448; // Line Descriptor
    2277: romdata_int <= 'h400;
    2278: romdata_int <= 'h1082;
    2279: romdata_int <= 'h4295;
    2280: romdata_int <= 'h448; // Line Descriptor
    2281: romdata_int <= 'h600;
    2282: romdata_int <= 'h76aa;
    2283: romdata_int <= 'h686c;
    2284: romdata_int <= 'h448; // Line Descriptor
    2285: romdata_int <= 'h800;
    2286: romdata_int <= 'hd1;
    2287: romdata_int <= 'h54b9;
    2288: romdata_int <= 'h448; // Line Descriptor
    2289: romdata_int <= 'ha00;
    2290: romdata_int <= 'h1900;
    2291: romdata_int <= 'h2156;
    2292: romdata_int <= 'h448; // Line Descriptor
    2293: romdata_int <= 'hc00;
    2294: romdata_int <= 'h4f20;
    2295: romdata_int <= 'h2f0a;
    2296: romdata_int <= 'h448; // Line Descriptor
    2297: romdata_int <= 'he00;
    2298: romdata_int <= 'h4507;
    2299: romdata_int <= 'h3698;
    2300: romdata_int <= 'h448; // Line Descriptor
    2301: romdata_int <= 'h1000;
    2302: romdata_int <= 'h24a;
    2303: romdata_int <= 'h4d15;
    2304: romdata_int <= 'h448; // Line Descriptor
    2305: romdata_int <= 'h1200;
    2306: romdata_int <= 'h809c;
    2307: romdata_int <= 'hf03;
    2308: romdata_int <= 'h448; // Line Descriptor
    2309: romdata_int <= 'h1400;
    2310: romdata_int <= 'h8cd0;
    2311: romdata_int <= 'h871e;
    2312: romdata_int <= 'h448; // Line Descriptor
    2313: romdata_int <= 'h1600;
    2314: romdata_int <= 'h3865;
    2315: romdata_int <= 'h4933;
    2316: romdata_int <= 'h448; // Line Descriptor
    2317: romdata_int <= 'h1800;
    2318: romdata_int <= 'h8b31;
    2319: romdata_int <= 'hac9;
    2320: romdata_int <= 'h448; // Line Descriptor
    2321: romdata_int <= 'h1a00;
    2322: romdata_int <= 'h529a;
    2323: romdata_int <= 'h2c0a;
    2324: romdata_int <= 'h448; // Line Descriptor
    2325: romdata_int <= 'h1c00;
    2326: romdata_int <= 'hcb8;
    2327: romdata_int <= 'h7abf;
    2328: romdata_int <= 'h448; // Line Descriptor
    2329: romdata_int <= 'h1e00;
    2330: romdata_int <= 'h150b;
    2331: romdata_int <= 'h32b8;
    2332: romdata_int <= 'h448; // Line Descriptor
    2333: romdata_int <= 'h2000;
    2334: romdata_int <= 'h3e54;
    2335: romdata_int <= 'h3525;
    2336: romdata_int <= 'h448; // Line Descriptor
    2337: romdata_int <= 'h2200;
    2338: romdata_int <= 'h3d3c;
    2339: romdata_int <= 'h8850;
    2340: romdata_int <= 'h448; // Line Descriptor
    2341: romdata_int <= 'h2400;
    2342: romdata_int <= 'h5f12;
    2343: romdata_int <= 'h8e3a;
    2344: romdata_int <= 'h448; // Line Descriptor
    2345: romdata_int <= 'h2600;
    2346: romdata_int <= 'h817;
    2347: romdata_int <= 'h5b0d;
    2348: romdata_int <= 'h448; // Line Descriptor
    2349: romdata_int <= 'h2800;
    2350: romdata_int <= 'h163d;
    2351: romdata_int <= 'h6232;
    2352: romdata_int <= 'h448; // Line Descriptor
    2353: romdata_int <= 'h2a00;
    2354: romdata_int <= 'h66b9;
    2355: romdata_int <= 'h767;
    2356: romdata_int <= 'h448; // Line Descriptor
    2357: romdata_int <= 'h2c00;
    2358: romdata_int <= 'h253c;
    2359: romdata_int <= 'h512e;
    2360: romdata_int <= 'h448; // Line Descriptor
    2361: romdata_int <= 'h2e00;
    2362: romdata_int <= 'h3a95;
    2363: romdata_int <= 'h26c4;
    2364: romdata_int <= 'h448; // Line Descriptor
    2365: romdata_int <= 'h3000;
    2366: romdata_int <= 'h1edf;
    2367: romdata_int <= 'h232c;
    2368: romdata_int <= 'h448; // Line Descriptor
    2369: romdata_int <= 'h3200;
    2370: romdata_int <= 'h7258;
    2371: romdata_int <= 'h6a33;
    2372: romdata_int <= 'h448; // Line Descriptor
    2373: romdata_int <= 'h3400;
    2374: romdata_int <= 'h2a08;
    2375: romdata_int <= 'h3115;
    2376: romdata_int <= 'h448; // Line Descriptor
    2377: romdata_int <= 'h3600;
    2378: romdata_int <= 'h6e4f;
    2379: romdata_int <= 'h2870;
    2380: romdata_int <= 'h448; // Line Descriptor
    2381: romdata_int <= 'h3800;
    2382: romdata_int <= 'h45e;
    2383: romdata_int <= 'h5884;
    2384: romdata_int <= 'h448; // Line Descriptor
    2385: romdata_int <= 'h3a00;
    2386: romdata_int <= 'h4a3b;
    2387: romdata_int <= 'h5cf3;
    2388: romdata_int <= 'h448; // Line Descriptor
    2389: romdata_int <= 'h3c00;
    2390: romdata_int <= 'h40bc;
    2391: romdata_int <= 'h7f39;
    2392: romdata_int <= 'h448; // Line Descriptor
    2393: romdata_int <= 'h3e00;
    2394: romdata_int <= 'h7418;
    2395: romdata_int <= 'h1240;
    2396: romdata_int <= 'h448; // Line Descriptor
    2397: romdata_int <= 'h4000;
    2398: romdata_int <= 'h6d42;
    2399: romdata_int <= 'h70a1;
    2400: romdata_int <= 'h448; // Line Descriptor
    2401: romdata_int <= 'h4200;
    2402: romdata_int <= 'h5710;
    2403: romdata_int <= 'h1c1c;
    2404: romdata_int <= 'h448; // Line Descriptor
    2405: romdata_int <= 'h4400;
    2406: romdata_int <= 'h82bc;
    2407: romdata_int <= 'h84ba;
    2408: romdata_int <= 'h448; // Line Descriptor
    2409: romdata_int <= 'h4600;
    2410: romdata_int <= 'h78be;
    2411: romdata_int <= 'h60f0;
    2412: romdata_int <= 'h448; // Line Descriptor
    2413: romdata_int <= 'h4800;
    2414: romdata_int <= 'h395b;
    2415: romdata_int <= 'h60c1;
    2416: romdata_int <= 'h448; // Line Descriptor
    2417: romdata_int <= 'h4a00;
    2418: romdata_int <= 'h6338;
    2419: romdata_int <= 'h7e5c;
    2420: romdata_int <= 'h448; // Line Descriptor
    2421: romdata_int <= 'h4c00;
    2422: romdata_int <= 'h4c44;
    2423: romdata_int <= 'h76ae;
    2424: romdata_int <= 'h448; // Line Descriptor
    2425: romdata_int <= 'h4e00;
    2426: romdata_int <= 'h3b26;
    2427: romdata_int <= 'h2a47;
    2428: romdata_int <= 'h448; // Line Descriptor
    2429: romdata_int <= 'h5000;
    2430: romdata_int <= 'h333b;
    2431: romdata_int <= 'h3460;
    2432: romdata_int <= 'h448; // Line Descriptor
    2433: romdata_int <= 'h5200;
    2434: romdata_int <= 'h5c68;
    2435: romdata_int <= 'h1356;
    2436: romdata_int <= 'h448; // Line Descriptor
    2437: romdata_int <= 'h5400;
    2438: romdata_int <= 'h8152;
    2439: romdata_int <= 'h6ab1;
    2440: romdata_int <= 'h448; // Line Descriptor
    2441: romdata_int <= 'h5600;
    2442: romdata_int <= 'h2f30;
    2443: romdata_int <= 'h1165;
    2444: romdata_int <= 'h448; // Line Descriptor
    2445: romdata_int <= 'h5800;
    2446: romdata_int <= 'h1ea7;
    2447: romdata_int <= 'h780f;
    2448: romdata_int <= 'h448; // Line Descriptor
    2449: romdata_int <= 'h5a00;
    2450: romdata_int <= 'h5551;
    2451: romdata_int <= 'h1a0e;
    2452: romdata_int <= 'h448; // Line Descriptor
    2453: romdata_int <= 'h5c00;
    2454: romdata_int <= 'h58c2;
    2455: romdata_int <= 'h1720;
    2456: romdata_int <= 'h448; // Line Descriptor
    2457: romdata_int <= 'h5e00;
    2458: romdata_int <= 'h429c;
    2459: romdata_int <= 'h36d3;
    2460: romdata_int <= 'h448; // Line Descriptor
    2461: romdata_int <= 'h6000;
    2462: romdata_int <= 'h7c40;
    2463: romdata_int <= 'h66d7;
    2464: romdata_int <= 'h448; // Line Descriptor
    2465: romdata_int <= 'h6200;
    2466: romdata_int <= 'h7282;
    2467: romdata_int <= 'h3ec7;
    2468: romdata_int <= 'h448; // Line Descriptor
    2469: romdata_int <= 'h6400;
    2470: romdata_int <= 'h4e21;
    2471: romdata_int <= 'h305a;
    2472: romdata_int <= 'h448; // Line Descriptor
    2473: romdata_int <= 'h6600;
    2474: romdata_int <= 'h695a;
    2475: romdata_int <= 'h8556;
    2476: romdata_int <= 'h448; // Line Descriptor
    2477: romdata_int <= 'h6800;
    2478: romdata_int <= 'h56c8;
    2479: romdata_int <= 'h407a;
    2480: romdata_int <= 'h448; // Line Descriptor
    2481: romdata_int <= 'h6a00;
    2482: romdata_int <= 'h1c60;
    2483: romdata_int <= 'h8611;
    2484: romdata_int <= 'h448; // Line Descriptor
    2485: romdata_int <= 'h6c00;
    2486: romdata_int <= 'h2256;
    2487: romdata_int <= 'h8d20;
    2488: romdata_int <= 'h448; // Line Descriptor
    2489: romdata_int <= 'h6e00;
    2490: romdata_int <= 'h26c1;
    2491: romdata_int <= 'h5e38;
    2492: romdata_int <= 'h448; // Line Descriptor
    2493: romdata_int <= 'h7000;
    2494: romdata_int <= 'h553;
    2495: romdata_int <= 'h28b7;
    2496: romdata_int <= 'h448; // Line Descriptor
    2497: romdata_int <= 'h7200;
    2498: romdata_int <= 'h52bb;
    2499: romdata_int <= 'h8a54;
    2500: romdata_int <= 'h448; // Line Descriptor
    2501: romdata_int <= 'h7400;
    2502: romdata_int <= 'ha89;
    2503: romdata_int <= 'h1872;
    2504: romdata_int <= 'h448; // Line Descriptor
    2505: romdata_int <= 'h7600;
    2506: romdata_int <= 'h7415;
    2507: romdata_int <= 'h8853;
    2508: romdata_int <= 'h448; // Line Descriptor
    2509: romdata_int <= 'h7800;
    2510: romdata_int <= 'h966;
    2511: romdata_int <= 'h46f1;
    2512: romdata_int <= 'h448; // Line Descriptor
    2513: romdata_int <= 'h7a00;
    2514: romdata_int <= 'hf1f;
    2515: romdata_int <= 'h35a;
    2516: romdata_int <= 'h448; // Line Descriptor
    2517: romdata_int <= 'h7c00;
    2518: romdata_int <= 'hd55;
    2519: romdata_int <= 'h8f1d;
    2520: romdata_int <= 'h448; // Line Descriptor
    2521: romdata_int <= 'h7e00;
    2522: romdata_int <= 'h24ac;
    2523: romdata_int <= 'h3c33;
    2524: romdata_int <= 'h448; // Line Descriptor
    2525: romdata_int <= 'h8000;
    2526: romdata_int <= 'h4473;
    2527: romdata_int <= 'h7a12;
    2528: romdata_int <= 'h448; // Line Descriptor
    2529: romdata_int <= 'h8200;
    2530: romdata_int <= 'h6f16;
    2531: romdata_int <= 'hcb;
    2532: romdata_int <= 'h448; // Line Descriptor
    2533: romdata_int <= 'h8400;
    2534: romdata_int <= 'h2cec;
    2535: romdata_int <= 'h2033;
    2536: romdata_int <= 'h448; // Line Descriptor
    2537: romdata_int <= 'h8600;
    2538: romdata_int <= 'h4b13;
    2539: romdata_int <= 'h140d;
    2540: romdata_int <= 'h448; // Line Descriptor
    2541: romdata_int <= 'h8800;
    2542: romdata_int <= 'h6d3;
    2543: romdata_int <= 'h50a8;
    2544: romdata_int <= 'h448; // Line Descriptor
    2545: romdata_int <= 'h8a00;
    2546: romdata_int <= 'h6c6b;
    2547: romdata_int <= 'h713c;
    2548: romdata_int <= 'h448; // Line Descriptor
    2549: romdata_int <= 'h8c00;
    2550: romdata_int <= 'h4831;
    2551: romdata_int <= 'h5a28;
    2552: romdata_int <= 'h548; // Line Descriptor
    2553: romdata_int <= 'h8e00;
    2554: romdata_int <= 'h642f;
    2555: romdata_int <= 'h826b;
    2556: romdata_int <= 'h183c; // Line Descriptor
    2557: romdata_int <= 'h0;
    2558: romdata_int <= 'h66ae;
    2559: romdata_int <= 'h2f0b;
    2560: romdata_int <= 'h3408;
    2561: romdata_int <= 'h5cd5;
    2562: romdata_int <= 'h3286;
    2563: romdata_int <= 'hc89;
    2564: romdata_int <= 'he2e;
    2565: romdata_int <= 'h4;
    2566: romdata_int <= 'h1b37;
    2567: romdata_int <= 'h4e9a;
    2568: romdata_int <= 'h26b0;
    2569: romdata_int <= 'h615c;
    2570: romdata_int <= 'h183c; // Line Descriptor
    2571: romdata_int <= 'h200;
    2572: romdata_int <= 'h7728;
    2573: romdata_int <= 'h428a;
    2574: romdata_int <= 'h1a6b;
    2575: romdata_int <= 'h5867;
    2576: romdata_int <= 'h2855;
    2577: romdata_int <= 'h861;
    2578: romdata_int <= 'h40d5;
    2579: romdata_int <= 'h371e;
    2580: romdata_int <= 'h50a5;
    2581: romdata_int <= 'hee0;
    2582: romdata_int <= 'h32e6;
    2583: romdata_int <= 'h734;
    2584: romdata_int <= 'h183c; // Line Descriptor
    2585: romdata_int <= 'h400;
    2586: romdata_int <= 'h232b;
    2587: romdata_int <= 'h3064;
    2588: romdata_int <= 'h5290;
    2589: romdata_int <= 'h3936;
    2590: romdata_int <= 'h1cd5;
    2591: romdata_int <= 'h4662;
    2592: romdata_int <= 'h70f2;
    2593: romdata_int <= 'h64b6;
    2594: romdata_int <= 'h8c9;
    2595: romdata_int <= 'h4b54;
    2596: romdata_int <= 'h1e4a;
    2597: romdata_int <= 'h1677;
    2598: romdata_int <= 'h183c; // Line Descriptor
    2599: romdata_int <= 'h600;
    2600: romdata_int <= 'h4b49;
    2601: romdata_int <= 'h667;
    2602: romdata_int <= 'h18a6;
    2603: romdata_int <= 'h20f2;
    2604: romdata_int <= 'h2c88;
    2605: romdata_int <= 'h6327;
    2606: romdata_int <= 'h2bd;
    2607: romdata_int <= 'h485c;
    2608: romdata_int <= 'h7648;
    2609: romdata_int <= 'h4522;
    2610: romdata_int <= 'h7301;
    2611: romdata_int <= 'h6934;
    2612: romdata_int <= 'h183c; // Line Descriptor
    2613: romdata_int <= 'h800;
    2614: romdata_int <= 'h3e4d;
    2615: romdata_int <= 'h1348;
    2616: romdata_int <= 'h601a;
    2617: romdata_int <= 'h760a;
    2618: romdata_int <= 'h3716;
    2619: romdata_int <= 'h6eee;
    2620: romdata_int <= 'h2e66;
    2621: romdata_int <= 'h7432;
    2622: romdata_int <= 'h4cf3;
    2623: romdata_int <= 'h1d2a;
    2624: romdata_int <= 'h5958;
    2625: romdata_int <= 'h3458;
    2626: romdata_int <= 'h183c; // Line Descriptor
    2627: romdata_int <= 'ha00;
    2628: romdata_int <= 'h74a2;
    2629: romdata_int <= 'h402a;
    2630: romdata_int <= 'h48c9;
    2631: romdata_int <= 'h12ce;
    2632: romdata_int <= 'h24fd;
    2633: romdata_int <= 'h3d19;
    2634: romdata_int <= 'h6650;
    2635: romdata_int <= 'h6233;
    2636: romdata_int <= 'h281c;
    2637: romdata_int <= 'hb38;
    2638: romdata_int <= 'h2221;
    2639: romdata_int <= 'h5508;
    2640: romdata_int <= 'h183c; // Line Descriptor
    2641: romdata_int <= 'hc00;
    2642: romdata_int <= 'hc08;
    2643: romdata_int <= 'h6665;
    2644: romdata_int <= 'h6e5;
    2645: romdata_int <= 'h22c0;
    2646: romdata_int <= 'h165d;
    2647: romdata_int <= 'h6a7b;
    2648: romdata_int <= 'h5efd;
    2649: romdata_int <= 'h5aeb;
    2650: romdata_int <= 'h5618;
    2651: romdata_int <= 'h5e40;
    2652: romdata_int <= 'h3f22;
    2653: romdata_int <= 'h14cf;
    2654: romdata_int <= 'h183c; // Line Descriptor
    2655: romdata_int <= 'he00;
    2656: romdata_int <= 'hf58;
    2657: romdata_int <= 'h3eee;
    2658: romdata_int <= 'h44c3;
    2659: romdata_int <= 'h5045;
    2660: romdata_int <= 'h1487;
    2661: romdata_int <= 'ha5c;
    2662: romdata_int <= 'h2aca;
    2663: romdata_int <= 'h5306;
    2664: romdata_int <= 'h337;
    2665: romdata_int <= 'h2b33;
    2666: romdata_int <= 'h12b0;
    2667: romdata_int <= 'h4088;
    2668: romdata_int <= 'h183c; // Line Descriptor
    2669: romdata_int <= 'h1000;
    2670: romdata_int <= 'h163f;
    2671: romdata_int <= 'h76f5;
    2672: romdata_int <= 'h30fe;
    2673: romdata_int <= 'h754b;
    2674: romdata_int <= 'h68a8;
    2675: romdata_int <= 'h497;
    2676: romdata_int <= 'h64a6;
    2677: romdata_int <= 'hcd5;
    2678: romdata_int <= 'h6eb1;
    2679: romdata_int <= 'h2ca1;
    2680: romdata_int <= 'h5d40;
    2681: romdata_int <= 'h6c5a;
    2682: romdata_int <= 'h183c; // Line Descriptor
    2683: romdata_int <= 'h1200;
    2684: romdata_int <= 'h3345;
    2685: romdata_int <= 'ha9e;
    2686: romdata_int <= 'h4a81;
    2687: romdata_int <= 'h274d;
    2688: romdata_int <= 'h4c8b;
    2689: romdata_int <= 'h3a99;
    2690: romdata_int <= 'h5634;
    2691: romdata_int <= 'h1951;
    2692: romdata_int <= 'h3c6f;
    2693: romdata_int <= 'h2513;
    2694: romdata_int <= 'h700b;
    2695: romdata_int <= 'h427a;
    2696: romdata_int <= 'h183c; // Line Descriptor
    2697: romdata_int <= 'h1400;
    2698: romdata_int <= 'h384c;
    2699: romdata_int <= 'h626f;
    2700: romdata_int <= 'h5550;
    2701: romdata_int <= 'h5ab5;
    2702: romdata_int <= 'h1e0f;
    2703: romdata_int <= 'h7247;
    2704: romdata_int <= 'h42b8;
    2705: romdata_int <= 'h20e2;
    2706: romdata_int <= 'h6b11;
    2707: romdata_int <= 'h1006;
    2708: romdata_int <= 'h383a;
    2709: romdata_int <= 'h6760;
    2710: romdata_int <= 'h183c; // Line Descriptor
    2711: romdata_int <= 'h1600;
    2712: romdata_int <= 'h40ea;
    2713: romdata_int <= 'h1a43;
    2714: romdata_int <= 'h4f4c;
    2715: romdata_int <= 'h10d2;
    2716: romdata_int <= 'h3e0a;
    2717: romdata_int <= 'h6d44;
    2718: romdata_int <= 'hec;
    2719: romdata_int <= 'h3a89;
    2720: romdata_int <= 'h2eaa;
    2721: romdata_int <= 'h3166;
    2722: romdata_int <= 'h46ce;
    2723: romdata_int <= 'h448;
    2724: romdata_int <= 'h43c; // Line Descriptor
    2725: romdata_int <= 'h1800;
    2726: romdata_int <= 'he6;
    2727: romdata_int <= 'h2ec;
    2728: romdata_int <= 'h43c; // Line Descriptor
    2729: romdata_int <= 'h1a00;
    2730: romdata_int <= 'h1031;
    2731: romdata_int <= 'h5ea0;
    2732: romdata_int <= 'h43c; // Line Descriptor
    2733: romdata_int <= 'h1c00;
    2734: romdata_int <= 'h6af4;
    2735: romdata_int <= 'hf0b;
    2736: romdata_int <= 'h43c; // Line Descriptor
    2737: romdata_int <= 'h1e00;
    2738: romdata_int <= 'h5d55;
    2739: romdata_int <= 'h54b8;
    2740: romdata_int <= 'h43c; // Line Descriptor
    2741: romdata_int <= 'h2000;
    2742: romdata_int <= 'h613;
    2743: romdata_int <= 'h2896;
    2744: romdata_int <= 'h43c; // Line Descriptor
    2745: romdata_int <= 'h2200;
    2746: romdata_int <= 'h2e1;
    2747: romdata_int <= 'h6c42;
    2748: romdata_int <= 'h43c; // Line Descriptor
    2749: romdata_int <= 'h2400;
    2750: romdata_int <= 'h6019;
    2751: romdata_int <= 'h3c24;
    2752: romdata_int <= 'h43c; // Line Descriptor
    2753: romdata_int <= 'h2600;
    2754: romdata_int <= 'h48cb;
    2755: romdata_int <= 'h2167;
    2756: romdata_int <= 'h43c; // Line Descriptor
    2757: romdata_int <= 'h2800;
    2758: romdata_int <= 'h6e22;
    2759: romdata_int <= 'h4b4b;
    2760: romdata_int <= 'h43c; // Line Descriptor
    2761: romdata_int <= 'h2a00;
    2762: romdata_int <= 'h6245;
    2763: romdata_int <= 'h4c84;
    2764: romdata_int <= 'h43c; // Line Descriptor
    2765: romdata_int <= 'h2c00;
    2766: romdata_int <= 'h5109;
    2767: romdata_int <= 'h38a7;
    2768: romdata_int <= 'h43c; // Line Descriptor
    2769: romdata_int <= 'h2e00;
    2770: romdata_int <= 'h4608;
    2771: romdata_int <= 'h1cd2;
    2772: romdata_int <= 'h43c; // Line Descriptor
    2773: romdata_int <= 'h3000;
    2774: romdata_int <= 'h528d;
    2775: romdata_int <= 'h648c;
    2776: romdata_int <= 'h43c; // Line Descriptor
    2777: romdata_int <= 'h3200;
    2778: romdata_int <= 'h1f25;
    2779: romdata_int <= 'h5917;
    2780: romdata_int <= 'h43c; // Line Descriptor
    2781: romdata_int <= 'h3400;
    2782: romdata_int <= 'h4262;
    2783: romdata_int <= 'h468d;
    2784: romdata_int <= 'h43c; // Line Descriptor
    2785: romdata_int <= 'h3600;
    2786: romdata_int <= 'h1d11;
    2787: romdata_int <= 'h56ad;
    2788: romdata_int <= 'h43c; // Line Descriptor
    2789: romdata_int <= 'h3800;
    2790: romdata_int <= 'h3a7b;
    2791: romdata_int <= 'h2a74;
    2792: romdata_int <= 'h43c; // Line Descriptor
    2793: romdata_int <= 'h3a00;
    2794: romdata_int <= 'h246f;
    2795: romdata_int <= 'h4f09;
    2796: romdata_int <= 'h43c; // Line Descriptor
    2797: romdata_int <= 'h3c00;
    2798: romdata_int <= 'h953;
    2799: romdata_int <= 'h36d8;
    2800: romdata_int <= 'h43c; // Line Descriptor
    2801: romdata_int <= 'h3e00;
    2802: romdata_int <= 'h6429;
    2803: romdata_int <= 'h10f3;
    2804: romdata_int <= 'h43c; // Line Descriptor
    2805: romdata_int <= 'h4000;
    2806: romdata_int <= 'h4d2a;
    2807: romdata_int <= 'h6e6e;
    2808: romdata_int <= 'h43c; // Line Descriptor
    2809: romdata_int <= 'h4200;
    2810: romdata_int <= 'h566f;
    2811: romdata_int <= 'h1744;
    2812: romdata_int <= 'h43c; // Line Descriptor
    2813: romdata_int <= 'h4400;
    2814: romdata_int <= 'h2008;
    2815: romdata_int <= 'h2246;
    2816: romdata_int <= 'h43c; // Line Descriptor
    2817: romdata_int <= 'h4600;
    2818: romdata_int <= 'h3c79;
    2819: romdata_int <= 'hc60;
    2820: romdata_int <= 'h43c; // Line Descriptor
    2821: romdata_int <= 'h4800;
    2822: romdata_int <= 'h2aaf;
    2823: romdata_int <= 'h5a94;
    2824: romdata_int <= 'h43c; // Line Descriptor
    2825: romdata_int <= 'h4a00;
    2826: romdata_int <= 'h4f53;
    2827: romdata_int <= 'h32c6;
    2828: romdata_int <= 'h43c; // Line Descriptor
    2829: romdata_int <= 'h4c00;
    2830: romdata_int <= 'h1444;
    2831: romdata_int <= 'h2461;
    2832: romdata_int <= 'h43c; // Line Descriptor
    2833: romdata_int <= 'h4e00;
    2834: romdata_int <= 'h53e;
    2835: romdata_int <= 'h11c;
    2836: romdata_int <= 'h43c; // Line Descriptor
    2837: romdata_int <= 'h5000;
    2838: romdata_int <= 'h1b51;
    2839: romdata_int <= 'h68cd;
    2840: romdata_int <= 'h43c; // Line Descriptor
    2841: romdata_int <= 'h5200;
    2842: romdata_int <= 'h5b42;
    2843: romdata_int <= 'h5d45;
    2844: romdata_int <= 'h43c; // Line Descriptor
    2845: romdata_int <= 'h5400;
    2846: romdata_int <= 'h1268;
    2847: romdata_int <= 'h153d;
    2848: romdata_int <= 'h43c; // Line Descriptor
    2849: romdata_int <= 'h5600;
    2850: romdata_int <= 'h72b7;
    2851: romdata_int <= 'h6b3f;
    2852: romdata_int <= 'h43c; // Line Descriptor
    2853: romdata_int <= 'h5800;
    2854: romdata_int <= 'h2949;
    2855: romdata_int <= 'h18c4;
    2856: romdata_int <= 'h43c; // Line Descriptor
    2857: romdata_int <= 'h5a00;
    2858: romdata_int <= 'h3147;
    2859: romdata_int <= 'h607b;
    2860: romdata_int <= 'h43c; // Line Descriptor
    2861: romdata_int <= 'h5c00;
    2862: romdata_int <= 'h710b;
    2863: romdata_int <= 'h523a;
    2864: romdata_int <= 'h43c; // Line Descriptor
    2865: romdata_int <= 'h5e00;
    2866: romdata_int <= 'h26c4;
    2867: romdata_int <= 'h55f;
    2868: romdata_int <= 'h43c; // Line Descriptor
    2869: romdata_int <= 'h6000;
    2870: romdata_int <= 'h54d9;
    2871: romdata_int <= 'h2ca1;
    2872: romdata_int <= 'h43c; // Line Descriptor
    2873: romdata_int <= 'h6200;
    2874: romdata_int <= 'h6c94;
    2875: romdata_int <= 'h7256;
    2876: romdata_int <= 'h43c; // Line Descriptor
    2877: romdata_int <= 'h6400;
    2878: romdata_int <= 'h5eb8;
    2879: romdata_int <= 'h2637;
    2880: romdata_int <= 'h43c; // Line Descriptor
    2881: romdata_int <= 'h6600;
    2882: romdata_int <= 'h693a;
    2883: romdata_int <= 'h4848;
    2884: romdata_int <= 'h43c; // Line Descriptor
    2885: romdata_int <= 'h6800;
    2886: romdata_int <= 'h4483;
    2887: romdata_int <= 'h7440;
    2888: romdata_int <= 'h43c; // Line Descriptor
    2889: romdata_int <= 'h6a00;
    2890: romdata_int <= 'h2e63;
    2891: romdata_int <= 'h5048;
    2892: romdata_int <= 'h43c; // Line Descriptor
    2893: romdata_int <= 'h6c00;
    2894: romdata_int <= 'h347a;
    2895: romdata_int <= 'h34c3;
    2896: romdata_int <= 'h43c; // Line Descriptor
    2897: romdata_int <= 'h6e00;
    2898: romdata_int <= 'h2c56;
    2899: romdata_int <= 'h3a5d;
    2900: romdata_int <= 'h43c; // Line Descriptor
    2901: romdata_int <= 'h7000;
    2902: romdata_int <= 'h1828;
    2903: romdata_int <= 'h1f20;
    2904: romdata_int <= 'h43c; // Line Descriptor
    2905: romdata_int <= 'h7200;
    2906: romdata_int <= 'haa4;
    2907: romdata_int <= 'h4555;
    2908: romdata_int <= 'h43c; // Line Descriptor
    2909: romdata_int <= 'h7400;
    2910: romdata_int <= 'h366f;
    2911: romdata_int <= 'h81f;
    2912: romdata_int <= 'h43c; // Line Descriptor
    2913: romdata_int <= 'h7600;
    2914: romdata_int <= 'h5956;
    2915: romdata_int <= 'h7056;
    2916: romdata_int <= 'h43c; // Line Descriptor
    2917: romdata_int <= 'h0;
    2918: romdata_int <= 'h5d2f;
    2919: romdata_int <= 'h5f1e;
    2920: romdata_int <= 'h43c; // Line Descriptor
    2921: romdata_int <= 'h200;
    2922: romdata_int <= 'h289c;
    2923: romdata_int <= 'h5c89;
    2924: romdata_int <= 'h43c; // Line Descriptor
    2925: romdata_int <= 'h400;
    2926: romdata_int <= 'h6a75;
    2927: romdata_int <= 'ha33;
    2928: romdata_int <= 'h43c; // Line Descriptor
    2929: romdata_int <= 'h600;
    2930: romdata_int <= 'h1930;
    2931: romdata_int <= 'h72df;
    2932: romdata_int <= 'h43c; // Line Descriptor
    2933: romdata_int <= 'h800;
    2934: romdata_int <= 'h5298;
    2935: romdata_int <= 'h5504;
    2936: romdata_int <= 'h43c; // Line Descriptor
    2937: romdata_int <= 'ha00;
    2938: romdata_int <= 'h44b2;
    2939: romdata_int <= 'h1aa9;
    2940: romdata_int <= 'h43c; // Line Descriptor
    2941: romdata_int <= 'hc00;
    2942: romdata_int <= 'hac1;
    2943: romdata_int <= 'h2497;
    2944: romdata_int <= 'h43c; // Line Descriptor
    2945: romdata_int <= 'he00;
    2946: romdata_int <= 'h2659;
    2947: romdata_int <= 'h749c;
    2948: romdata_int <= 'h43c; // Line Descriptor
    2949: romdata_int <= 'h1000;
    2950: romdata_int <= 'h3096;
    2951: romdata_int <= 'h469e;
    2952: romdata_int <= 'h43c; // Line Descriptor
    2953: romdata_int <= 'h1200;
    2954: romdata_int <= 'hc14;
    2955: romdata_int <= 'h4510;
    2956: romdata_int <= 'h43c; // Line Descriptor
    2957: romdata_int <= 'h1400;
    2958: romdata_int <= 'h6cf9;
    2959: romdata_int <= 'h2c12;
    2960: romdata_int <= 'h43c; // Line Descriptor
    2961: romdata_int <= 'h1600;
    2962: romdata_int <= 'h1e9c;
    2963: romdata_int <= 'h495a;
    2964: romdata_int <= 'h43c; // Line Descriptor
    2965: romdata_int <= 'h1800;
    2966: romdata_int <= 'h90a;
    2967: romdata_int <= 'h3664;
    2968: romdata_int <= 'h43c; // Line Descriptor
    2969: romdata_int <= 'h1a00;
    2970: romdata_int <= 'h3af6;
    2971: romdata_int <= 'h406b;
    2972: romdata_int <= 'h43c; // Line Descriptor
    2973: romdata_int <= 'h1c00;
    2974: romdata_int <= 'h2c85;
    2975: romdata_int <= 'h6735;
    2976: romdata_int <= 'h43c; // Line Descriptor
    2977: romdata_int <= 'h1e00;
    2978: romdata_int <= 'h54f5;
    2979: romdata_int <= 'h62ea;
    2980: romdata_int <= 'h43c; // Line Descriptor
    2981: romdata_int <= 'h2000;
    2982: romdata_int <= 'h1a04;
    2983: romdata_int <= 'h5a32;
    2984: romdata_int <= 'h43c; // Line Descriptor
    2985: romdata_int <= 'h2200;
    2986: romdata_int <= 'h1c15;
    2987: romdata_int <= 'h3541;
    2988: romdata_int <= 'h43c; // Line Descriptor
    2989: romdata_int <= 'h2400;
    2990: romdata_int <= 'h22f6;
    2991: romdata_int <= 'h822;
    2992: romdata_int <= 'h43c; // Line Descriptor
    2993: romdata_int <= 'h2600;
    2994: romdata_int <= 'he8;
    2995: romdata_int <= 'ha5;
    2996: romdata_int <= 'h43c; // Line Descriptor
    2997: romdata_int <= 'h2800;
    2998: romdata_int <= 'h4007;
    2999: romdata_int <= 'h6c7a;
    3000: romdata_int <= 'h43c; // Line Descriptor
    3001: romdata_int <= 'h2a00;
    3002: romdata_int <= 'h352f;
    3003: romdata_int <= 'h2aa5;
    3004: romdata_int <= 'h43c; // Line Descriptor
    3005: romdata_int <= 'h2c00;
    3006: romdata_int <= 'h1666;
    3007: romdata_int <= 'h1c5a;
    3008: romdata_int <= 'h43c; // Line Descriptor
    3009: romdata_int <= 'h2e00;
    3010: romdata_int <= 'h72a7;
    3011: romdata_int <= 'hca2;
    3012: romdata_int <= 'h43c; // Line Descriptor
    3013: romdata_int <= 'h3000;
    3014: romdata_int <= 'h5ac8;
    3015: romdata_int <= 'h265b;
    3016: romdata_int <= 'h43c; // Line Descriptor
    3017: romdata_int <= 'h3200;
    3018: romdata_int <= 'h448;
    3019: romdata_int <= 'h1485;
    3020: romdata_int <= 'h43c; // Line Descriptor
    3021: romdata_int <= 'h3400;
    3022: romdata_int <= 'h2104;
    3023: romdata_int <= 'h3c5c;
    3024: romdata_int <= 'h43c; // Line Descriptor
    3025: romdata_int <= 'h3600;
    3026: romdata_int <= 'h2b03;
    3027: romdata_int <= 'h52b1;
    3028: romdata_int <= 'h43c; // Line Descriptor
    3029: romdata_int <= 'h3800;
    3030: romdata_int <= 'h2559;
    3031: romdata_int <= 'he7b;
    3032: romdata_int <= 'h43c; // Line Descriptor
    3033: romdata_int <= 'h3a00;
    3034: romdata_int <= 'h7429;
    3035: romdata_int <= 'h3139;
    3036: romdata_int <= 'h43c; // Line Descriptor
    3037: romdata_int <= 'h3c00;
    3038: romdata_int <= 'h5895;
    3039: romdata_int <= 'h282b;
    3040: romdata_int <= 'h43c; // Line Descriptor
    3041: romdata_int <= 'h3e00;
    3042: romdata_int <= 'h486c;
    3043: romdata_int <= 'h3b2a;
    3044: romdata_int <= 'h43c; // Line Descriptor
    3045: romdata_int <= 'h4000;
    3046: romdata_int <= 'h60b9;
    3047: romdata_int <= 'h4c01;
    3048: romdata_int <= 'h43c; // Line Descriptor
    3049: romdata_int <= 'h4200;
    3050: romdata_int <= 'h4f56;
    3051: romdata_int <= 'h583d;
    3052: romdata_int <= 'h43c; // Line Descriptor
    3053: romdata_int <= 'h4400;
    3054: romdata_int <= 'h147d;
    3055: romdata_int <= 'h121a;
    3056: romdata_int <= 'h43c; // Line Descriptor
    3057: romdata_int <= 'h4600;
    3058: romdata_int <= 'h510a;
    3059: romdata_int <= 'h68c2;
    3060: romdata_int <= 'h43c; // Line Descriptor
    3061: romdata_int <= 'h4800;
    3062: romdata_int <= 'h3698;
    3063: romdata_int <= 'h56ab;
    3064: romdata_int <= 'h43c; // Line Descriptor
    3065: romdata_int <= 'h4a00;
    3066: romdata_int <= 'h3d15;
    3067: romdata_int <= 'h1603;
    3068: romdata_int <= 'h43c; // Line Descriptor
    3069: romdata_int <= 'h4c00;
    3070: romdata_int <= 'h4b03;
    3071: romdata_int <= 'h3337;
    3072: romdata_int <= 'h43c; // Line Descriptor
    3073: romdata_int <= 'h4e00;
    3074: romdata_int <= 'hf1e;
    3075: romdata_int <= 'h4b5c;
    3076: romdata_int <= 'h43c; // Line Descriptor
    3077: romdata_int <= 'h5000;
    3078: romdata_int <= 'h7046;
    3079: romdata_int <= 'h3e38;
    3080: romdata_int <= 'h43c; // Line Descriptor
    3081: romdata_int <= 'h5200;
    3082: romdata_int <= 'h694e;
    3083: romdata_int <= 'h771e;
    3084: romdata_int <= 'h43c; // Line Descriptor
    3085: romdata_int <= 'h5400;
    3086: romdata_int <= 'h4c99;
    3087: romdata_int <= 'h2054;
    3088: romdata_int <= 'h43c; // Line Descriptor
    3089: romdata_int <= 'h5600;
    3090: romdata_int <= 'h1333;
    3091: romdata_int <= 'h188d;
    3092: romdata_int <= 'h43c; // Line Descriptor
    3093: romdata_int <= 'h5800;
    3094: romdata_int <= 'h42c9;
    3095: romdata_int <= 'h6b59;
    3096: romdata_int <= 'h43c; // Line Descriptor
    3097: romdata_int <= 'h5a00;
    3098: romdata_int <= 'h3310;
    3099: romdata_int <= 'h38d4;
    3100: romdata_int <= 'h43c; // Line Descriptor
    3101: romdata_int <= 'h5c00;
    3102: romdata_int <= 'h70b;
    3103: romdata_int <= 'h6eb8;
    3104: romdata_int <= 'h43c; // Line Descriptor
    3105: romdata_int <= 'h5e00;
    3106: romdata_int <= 'h1054;
    3107: romdata_int <= 'h1f25;
    3108: romdata_int <= 'h43c; // Line Descriptor
    3109: romdata_int <= 'h6000;
    3110: romdata_int <= 'h473c;
    3111: romdata_int <= 'h2250;
    3112: romdata_int <= 'h43c; // Line Descriptor
    3113: romdata_int <= 'h6200;
    3114: romdata_int <= 'h5712;
    3115: romdata_int <= 'h703a;
    3116: romdata_int <= 'h43c; // Line Descriptor
    3117: romdata_int <= 'h6400;
    3118: romdata_int <= 'h7617;
    3119: romdata_int <= 'h110d;
    3120: romdata_int <= 'h43c; // Line Descriptor
    3121: romdata_int <= 'h6600;
    3122: romdata_int <= 'h23d;
    3123: romdata_int <= 'h4e32;
    3124: romdata_int <= 'h43c; // Line Descriptor
    3125: romdata_int <= 'h6800;
    3126: romdata_int <= 'h653c;
    3127: romdata_int <= 'h32e;
    3128: romdata_int <= 'h43c; // Line Descriptor
    3129: romdata_int <= 'h6a00;
    3130: romdata_int <= 'h3895;
    3131: romdata_int <= 'h42c4;
    3132: romdata_int <= 'h43c; // Line Descriptor
    3133: romdata_int <= 'h6c00;
    3134: romdata_int <= 'h5edf;
    3135: romdata_int <= 'h72c;
    3136: romdata_int <= 'h43c; // Line Descriptor
    3137: romdata_int <= 'h6e00;
    3138: romdata_int <= 'h2e58;
    3139: romdata_int <= 'h2e33;
    3140: romdata_int <= 'h43c; // Line Descriptor
    3141: romdata_int <= 'h7000;
    3142: romdata_int <= 'h6608;
    3143: romdata_int <= 'h6115;
    3144: romdata_int <= 'h43c; // Line Descriptor
    3145: romdata_int <= 'h7200;
    3146: romdata_int <= 'h3e4f;
    3147: romdata_int <= 'h470;
    3148: romdata_int <= 'h43c; // Line Descriptor
    3149: romdata_int <= 'h7400;
    3150: romdata_int <= 'h6e5e;
    3151: romdata_int <= 'h5084;
    3152: romdata_int <= 'h53c; // Line Descriptor
    3153: romdata_int <= 'h7600;
    3154: romdata_int <= 'h623b;
    3155: romdata_int <= 'h64f3;
    3156: romdata_int <= 'h162d; // Line Descriptor
    3157: romdata_int <= 'h0;
    3158: romdata_int <= 'h508d;
    3159: romdata_int <= 'h34af;
    3160: romdata_int <= 'h3f44;
    3161: romdata_int <= 'h3129;
    3162: romdata_int <= 'h50f8;
    3163: romdata_int <= 'h1848;
    3164: romdata_int <= 'h2e74;
    3165: romdata_int <= 'h3a37;
    3166: romdata_int <= 'h2c3c;
    3167: romdata_int <= 'h1612;
    3168: romdata_int <= 'h4ea3;
    3169: romdata_int <= 'h162d; // Line Descriptor
    3170: romdata_int <= 'h200;
    3171: romdata_int <= 'h26fc;
    3172: romdata_int <= 'h563b;
    3173: romdata_int <= 'h5407;
    3174: romdata_int <= 'h1333;
    3175: romdata_int <= 'h4b1b;
    3176: romdata_int <= 'h58a0;
    3177: romdata_int <= 'h496;
    3178: romdata_int <= 'h1554;
    3179: romdata_int <= 'h5412;
    3180: romdata_int <= 'h2a2c;
    3181: romdata_int <= 'h40fd;
    3182: romdata_int <= 'h162d; // Line Descriptor
    3183: romdata_int <= 'h400;
    3184: romdata_int <= 'h40ae;
    3185: romdata_int <= 'h18b1;
    3186: romdata_int <= 'h2a8c;
    3187: romdata_int <= 'h2d2e;
    3188: romdata_int <= 'h50f;
    3189: romdata_int <= 'h941;
    3190: romdata_int <= 'h2350;
    3191: romdata_int <= 'h134;
    3192: romdata_int <= 'h5625;
    3193: romdata_int <= 'h128e;
    3194: romdata_int <= 'h452a;
    3195: romdata_int <= 'h162d; // Line Descriptor
    3196: romdata_int <= 'h600;
    3197: romdata_int <= 'h3c22;
    3198: romdata_int <= 'h1d06;
    3199: romdata_int <= 'h9b;
    3200: romdata_int <= 'h2327;
    3201: romdata_int <= 'h251;
    3202: romdata_int <= 'h4054;
    3203: romdata_int <= 'h54c2;
    3204: romdata_int <= 'h20a2;
    3205: romdata_int <= 'h4680;
    3206: romdata_int <= 'h233e;
    3207: romdata_int <= 'h48ae;
    3208: romdata_int <= 'h162d; // Line Descriptor
    3209: romdata_int <= 'h800;
    3210: romdata_int <= 'h2aa9;
    3211: romdata_int <= 'h2cfd;
    3212: romdata_int <= 'h2744;
    3213: romdata_int <= 'h1cd7;
    3214: romdata_int <= 'h1024;
    3215: romdata_int <= 'h562e;
    3216: romdata_int <= 'h12f0;
    3217: romdata_int <= 'h1ace;
    3218: romdata_int <= 'h1e1b;
    3219: romdata_int <= 'h3f52;
    3220: romdata_int <= 'h146c;
    3221: romdata_int <= 'h162d; // Line Descriptor
    3222: romdata_int <= 'ha00;
    3223: romdata_int <= 'h4623;
    3224: romdata_int <= 'h3a7e;
    3225: romdata_int <= 'h4960;
    3226: romdata_int <= 'h52d1;
    3227: romdata_int <= 'hb16;
    3228: romdata_int <= 'ha1f;
    3229: romdata_int <= 'h68c;
    3230: romdata_int <= 'h1678;
    3231: romdata_int <= 'hd3b;
    3232: romdata_int <= 'h2935;
    3233: romdata_int <= 'h2ea3;
    3234: romdata_int <= 'h162d; // Line Descriptor
    3235: romdata_int <= 'hc00;
    3236: romdata_int <= 'h125a;
    3237: romdata_int <= 'h20c4;
    3238: romdata_int <= 'h3c4b;
    3239: romdata_int <= 'h2eae;
    3240: romdata_int <= 'h36b1;
    3241: romdata_int <= 'h4954;
    3242: romdata_int <= 'h3c84;
    3243: romdata_int <= 'h24e6;
    3244: romdata_int <= 'h24e4;
    3245: romdata_int <= 'hd7;
    3246: romdata_int <= 'h2067;
    3247: romdata_int <= 'h162d; // Line Descriptor
    3248: romdata_int <= 'he00;
    3249: romdata_int <= 'h3e62;
    3250: romdata_int <= 'h658;
    3251: romdata_int <= 'h24cb;
    3252: romdata_int <= 'h4e2e;
    3253: romdata_int <= 'h4d19;
    3254: romdata_int <= 'h44a5;
    3255: romdata_int <= 'h1f0b;
    3256: romdata_int <= 'h350f;
    3257: romdata_int <= 'h580d;
    3258: romdata_int <= 'h552;
    3259: romdata_int <= 'h209;
    3260: romdata_int <= 'h162d; // Line Descriptor
    3261: romdata_int <= 'h1000;
    3262: romdata_int <= 'h2c85;
    3263: romdata_int <= 'h52ba;
    3264: romdata_int <= 'h1680;
    3265: romdata_int <= 'h404d;
    3266: romdata_int <= 'h60c;
    3267: romdata_int <= 'h373b;
    3268: romdata_int <= 'h2813;
    3269: romdata_int <= 'hccc;
    3270: romdata_int <= 'h328a;
    3271: romdata_int <= 'h735;
    3272: romdata_int <= 'h104f;
    3273: romdata_int <= 'h162d; // Line Descriptor
    3274: romdata_int <= 'h1200;
    3275: romdata_int <= 'h4a47;
    3276: romdata_int <= 'h1493;
    3277: romdata_int <= 'h326a;
    3278: romdata_int <= 'hc0c;
    3279: romdata_int <= 'h20d9;
    3280: romdata_int <= 'h22e;
    3281: romdata_int <= 'h2ca2;
    3282: romdata_int <= 'h304b;
    3283: romdata_int <= 'haa1;
    3284: romdata_int <= 'h366d;
    3285: romdata_int <= 'hf19;
    3286: romdata_int <= 'h162d; // Line Descriptor
    3287: romdata_int <= 'h1400;
    3288: romdata_int <= 'hc4;
    3289: romdata_int <= 'h10e0;
    3290: romdata_int <= 'h28f6;
    3291: romdata_int <= 'h89d;
    3292: romdata_int <= 'h1e92;
    3293: romdata_int <= 'h4f23;
    3294: romdata_int <= 'h42e1;
    3295: romdata_int <= 'h389f;
    3296: romdata_int <= 'h4c0a;
    3297: romdata_int <= 'h3ca5;
    3298: romdata_int <= 'h1acd;
    3299: romdata_int <= 'h162d; // Line Descriptor
    3300: romdata_int <= 'h1600;
    3301: romdata_int <= 'h1a2a;
    3302: romdata_int <= 'h24f0;
    3303: romdata_int <= 'h3a02;
    3304: romdata_int <= 'h4604;
    3305: romdata_int <= 'h56a7;
    3306: romdata_int <= 'h2af5;
    3307: romdata_int <= 'h50eb;
    3308: romdata_int <= 'h3300;
    3309: romdata_int <= 'h3148;
    3310: romdata_int <= 'h52b0;
    3311: romdata_int <= 'h95b;
    3312: romdata_int <= 'h162d; // Line Descriptor
    3313: romdata_int <= 'h1800;
    3314: romdata_int <= 'h1451;
    3315: romdata_int <= 'hcc2;
    3316: romdata_int <= 'h186d;
    3317: romdata_int <= 'h4560;
    3318: romdata_int <= 'h5871;
    3319: romdata_int <= 'h262f;
    3320: romdata_int <= 'h1d62;
    3321: romdata_int <= 'h1148;
    3322: romdata_int <= 'h509e;
    3323: romdata_int <= 'h4a3b;
    3324: romdata_int <= 'h3a20;
    3325: romdata_int <= 'h162d; // Line Descriptor
    3326: romdata_int <= 'h1a00;
    3327: romdata_int <= 'h48b8;
    3328: romdata_int <= 'h5054;
    3329: romdata_int <= 'h140b;
    3330: romdata_int <= 'h1ac6;
    3331: romdata_int <= 'he96;
    3332: romdata_int <= 'h5211;
    3333: romdata_int <= 'h4ab0;
    3334: romdata_int <= 'h3e5d;
    3335: romdata_int <= 'h275a;
    3336: romdata_int <= 'h1d26;
    3337: romdata_int <= 'h183a;
    3338: romdata_int <= 'h162d; // Line Descriptor
    3339: romdata_int <= 'h1c00;
    3340: romdata_int <= 'h2541;
    3341: romdata_int <= 'h4a6b;
    3342: romdata_int <= 'h395d;
    3343: romdata_int <= 'h3443;
    3344: romdata_int <= 'h42f8;
    3345: romdata_int <= 'h471d;
    3346: romdata_int <= 'h4d2f;
    3347: romdata_int <= 'heb5;
    3348: romdata_int <= 'h3491;
    3349: romdata_int <= 'h434f;
    3350: romdata_int <= 'h38c2;
    3351: romdata_int <= 'h42d; // Line Descriptor
    3352: romdata_int <= 'h1e00;
    3353: romdata_int <= 'h5845;
    3354: romdata_int <= 'h170a;
    3355: romdata_int <= 'h42d; // Line Descriptor
    3356: romdata_int <= 'h2000;
    3357: romdata_int <= 'hd2a;
    3358: romdata_int <= 'h2a99;
    3359: romdata_int <= 'h42d; // Line Descriptor
    3360: romdata_int <= 'h2200;
    3361: romdata_int <= 'h723;
    3362: romdata_int <= 'h4128;
    3363: romdata_int <= 'h42d; // Line Descriptor
    3364: romdata_int <= 'h2400;
    3365: romdata_int <= 'h3a2c;
    3366: romdata_int <= 'h1f41;
    3367: romdata_int <= 'h42d; // Line Descriptor
    3368: romdata_int <= 'h2600;
    3369: romdata_int <= 'hea0;
    3370: romdata_int <= 'h4e5f;
    3371: romdata_int <= 'h42d; // Line Descriptor
    3372: romdata_int <= 'h2800;
    3373: romdata_int <= 'h3649;
    3374: romdata_int <= 'h3c57;
    3375: romdata_int <= 'h42d; // Line Descriptor
    3376: romdata_int <= 'h2a00;
    3377: romdata_int <= 'h1062;
    3378: romdata_int <= 'h4c8a;
    3379: romdata_int <= 'h42d; // Line Descriptor
    3380: romdata_int <= 'h2c00;
    3381: romdata_int <= 'h1c3b;
    3382: romdata_int <= 'h3336;
    3383: romdata_int <= 'h42d; // Line Descriptor
    3384: romdata_int <= 'h2e00;
    3385: romdata_int <= 'h16a8;
    3386: romdata_int <= 'h2ec8;
    3387: romdata_int <= 'h42d; // Line Descriptor
    3388: romdata_int <= 'h3000;
    3389: romdata_int <= 'h553a;
    3390: romdata_int <= 'h5441;
    3391: romdata_int <= 'h42d; // Line Descriptor
    3392: romdata_int <= 'h3200;
    3393: romdata_int <= 'h34a1;
    3394: romdata_int <= 'h389e;
    3395: romdata_int <= 'h42d; // Line Descriptor
    3396: romdata_int <= 'h3400;
    3397: romdata_int <= 'h1e88;
    3398: romdata_int <= 'h472f;
    3399: romdata_int <= 'h42d; // Line Descriptor
    3400: romdata_int <= 'h3600;
    3401: romdata_int <= 'h28a6;
    3402: romdata_int <= 'h3143;
    3403: romdata_int <= 'h42d; // Line Descriptor
    3404: romdata_int <= 'h3800;
    3405: romdata_int <= 'h22c0;
    3406: romdata_int <= 'h4836;
    3407: romdata_int <= 'h42d; // Line Descriptor
    3408: romdata_int <= 'h3a00;
    3409: romdata_int <= 'h8bf;
    3410: romdata_int <= 'h131d;
    3411: romdata_int <= 'h42d; // Line Descriptor
    3412: romdata_int <= 'h3c00;
    3413: romdata_int <= 'ha4d;
    3414: romdata_int <= 'h446;
    3415: romdata_int <= 'h42d; // Line Descriptor
    3416: romdata_int <= 'h3e00;
    3417: romdata_int <= 'h1935;
    3418: romdata_int <= 'h61;
    3419: romdata_int <= 'h42d; // Line Descriptor
    3420: romdata_int <= 'h4000;
    3421: romdata_int <= 'h4e85;
    3422: romdata_int <= 'hb31;
    3423: romdata_int <= 'h42d; // Line Descriptor
    3424: romdata_int <= 'h4200;
    3425: romdata_int <= 'h4cf3;
    3426: romdata_int <= 'hf3b;
    3427: romdata_int <= 'h42d; // Line Descriptor
    3428: romdata_int <= 'h4400;
    3429: romdata_int <= 'h4436;
    3430: romdata_int <= 'h3724;
    3431: romdata_int <= 'h42d; // Line Descriptor
    3432: romdata_int <= 'h4600;
    3433: romdata_int <= 'h2075;
    3434: romdata_int <= 'h274e;
    3435: romdata_int <= 'h42d; // Line Descriptor
    3436: romdata_int <= 'h4800;
    3437: romdata_int <= 'h2e18;
    3438: romdata_int <= 'h829;
    3439: romdata_int <= 'h42d; // Line Descriptor
    3440: romdata_int <= 'h4a00;
    3441: romdata_int <= 'h422d;
    3442: romdata_int <= 'h4417;
    3443: romdata_int <= 'h42d; // Line Descriptor
    3444: romdata_int <= 'h4c00;
    3445: romdata_int <= 'h30d6;
    3446: romdata_int <= 'h2887;
    3447: romdata_int <= 'h42d; // Line Descriptor
    3448: romdata_int <= 'h4e00;
    3449: romdata_int <= 'h33e;
    3450: romdata_int <= 'h22aa;
    3451: romdata_int <= 'h42d; // Line Descriptor
    3452: romdata_int <= 'h5000;
    3453: romdata_int <= 'h55b;
    3454: romdata_int <= 'h2b5;
    3455: romdata_int <= 'h42d; // Line Descriptor
    3456: romdata_int <= 'h5200;
    3457: romdata_int <= 'h5665;
    3458: romdata_int <= 'h1af9;
    3459: romdata_int <= 'h42d; // Line Descriptor
    3460: romdata_int <= 'h5400;
    3461: romdata_int <= 'h332f;
    3462: romdata_int <= 'h428a;
    3463: romdata_int <= 'h42d; // Line Descriptor
    3464: romdata_int <= 'h5600;
    3465: romdata_int <= 'h38be;
    3466: romdata_int <= 'h58ae;
    3467: romdata_int <= 'h42d; // Line Descriptor
    3468: romdata_int <= 'h5800;
    3469: romdata_int <= 'h5304;
    3470: romdata_int <= 'h3e3b;
    3471: romdata_int <= 'h42d; // Line Descriptor
    3472: romdata_int <= 'h0;
    3473: romdata_int <= 'h4016;
    3474: romdata_int <= 'h81c;
    3475: romdata_int <= 'h42d; // Line Descriptor
    3476: romdata_int <= 'h200;
    3477: romdata_int <= 'h918;
    3478: romdata_int <= 'h28dd;
    3479: romdata_int <= 'h42d; // Line Descriptor
    3480: romdata_int <= 'h400;
    3481: romdata_int <= 'h36b6;
    3482: romdata_int <= 'he3c;
    3483: romdata_int <= 'h42d; // Line Descriptor
    3484: romdata_int <= 'h600;
    3485: romdata_int <= 'hc46;
    3486: romdata_int <= 'h706;
    3487: romdata_int <= 'h42d; // Line Descriptor
    3488: romdata_int <= 'h800;
    3489: romdata_int <= 'h4e07;
    3490: romdata_int <= 'h3a21;
    3491: romdata_int <= 'h42d; // Line Descriptor
    3492: romdata_int <= 'ha00;
    3493: romdata_int <= 'h69b;
    3494: romdata_int <= 'h2538;
    3495: romdata_int <= 'h42d; // Line Descriptor
    3496: romdata_int <= 'hc00;
    3497: romdata_int <= 'h4b0;
    3498: romdata_int <= 'h1d65;
    3499: romdata_int <= 'h42d; // Line Descriptor
    3500: romdata_int <= 'he00;
    3501: romdata_int <= 'h194f;
    3502: romdata_int <= 'h430d;
    3503: romdata_int <= 'h42d; // Line Descriptor
    3504: romdata_int <= 'h1000;
    3505: romdata_int <= 'h1a70;
    3506: romdata_int <= 'h468f;
    3507: romdata_int <= 'h42d; // Line Descriptor
    3508: romdata_int <= 'h1200;
    3509: romdata_int <= 'h5519;
    3510: romdata_int <= 'h4b4b;
    3511: romdata_int <= 'h42d; // Line Descriptor
    3512: romdata_int <= 'h1400;
    3513: romdata_int <= 'h2f57;
    3514: romdata_int <= 'h1027;
    3515: romdata_int <= 'h42d; // Line Descriptor
    3516: romdata_int <= 'h1600;
    3517: romdata_int <= 'h2ab4;
    3518: romdata_int <= 'h1626;
    3519: romdata_int <= 'h42d; // Line Descriptor
    3520: romdata_int <= 'h1800;
    3521: romdata_int <= 'h1714;
    3522: romdata_int <= 'h120c;
    3523: romdata_int <= 'h42d; // Line Descriptor
    3524: romdata_int <= 'h1a00;
    3525: romdata_int <= 'h445b;
    3526: romdata_int <= 'h349d;
    3527: romdata_int <= 'h42d; // Line Descriptor
    3528: romdata_int <= 'h1c00;
    3529: romdata_int <= 'h3e1f;
    3530: romdata_int <= 'hbb;
    3531: romdata_int <= 'h42d; // Line Descriptor
    3532: romdata_int <= 'h1e00;
    3533: romdata_int <= 'h24d9;
    3534: romdata_int <= 'h58a8;
    3535: romdata_int <= 'h42d; // Line Descriptor
    3536: romdata_int <= 'h2000;
    3537: romdata_int <= 'h508b;
    3538: romdata_int <= 'h44fb;
    3539: romdata_int <= 'h42d; // Line Descriptor
    3540: romdata_int <= 'h2200;
    3541: romdata_int <= 'h1c1f;
    3542: romdata_int <= 'h30c;
    3543: romdata_int <= 'h42d; // Line Descriptor
    3544: romdata_int <= 'h2400;
    3545: romdata_int <= 'h14b3;
    3546: romdata_int <= 'h54c9;
    3547: romdata_int <= 'h42d; // Line Descriptor
    3548: romdata_int <= 'h2600;
    3549: romdata_int <= 'h4c40;
    3550: romdata_int <= 'h2ebb;
    3551: romdata_int <= 'h42d; // Line Descriptor
    3552: romdata_int <= 'h2800;
    3553: romdata_int <= 'h421c;
    3554: romdata_int <= 'h3d39;
    3555: romdata_int <= 'h42d; // Line Descriptor
    3556: romdata_int <= 'h2a00;
    3557: romdata_int <= 'he57;
    3558: romdata_int <= 'h4933;
    3559: romdata_int <= 'h42d; // Line Descriptor
    3560: romdata_int <= 'h2c00;
    3561: romdata_int <= 'h3455;
    3562: romdata_int <= 'h5058;
    3563: romdata_int <= 'h42d; // Line Descriptor
    3564: romdata_int <= 'h2e00;
    3565: romdata_int <= 'h1e82;
    3566: romdata_int <= 'h1a27;
    3567: romdata_int <= 'h42d; // Line Descriptor
    3568: romdata_int <= 'h3000;
    3569: romdata_int <= 'h3b;
    3570: romdata_int <= 'h234c;
    3571: romdata_int <= 'h42d; // Line Descriptor
    3572: romdata_int <= 'h3200;
    3573: romdata_int <= 'h3c7b;
    3574: romdata_int <= 'h408c;
    3575: romdata_int <= 'h42d; // Line Descriptor
    3576: romdata_int <= 'h3400;
    3577: romdata_int <= 'h385f;
    3578: romdata_int <= 'h3f18;
    3579: romdata_int <= 'h42d; // Line Descriptor
    3580: romdata_int <= 'h3600;
    3581: romdata_int <= 'h5702;
    3582: romdata_int <= 'h530f;
    3583: romdata_int <= 'h42d; // Line Descriptor
    3584: romdata_int <= 'h3800;
    3585: romdata_int <= 'hb64;
    3586: romdata_int <= 'h36a9;
    3587: romdata_int <= 'h42d; // Line Descriptor
    3588: romdata_int <= 'h3a00;
    3589: romdata_int <= 'h2867;
    3590: romdata_int <= 'h5739;
    3591: romdata_int <= 'h42d; // Line Descriptor
    3592: romdata_int <= 'h3c00;
    3593: romdata_int <= 'h58d4;
    3594: romdata_int <= 'h3923;
    3595: romdata_int <= 'h42d; // Line Descriptor
    3596: romdata_int <= 'h3e00;
    3597: romdata_int <= 'h4b36;
    3598: romdata_int <= 'h18d5;
    3599: romdata_int <= 'h42d; // Line Descriptor
    3600: romdata_int <= 'h4000;
    3601: romdata_int <= 'h2756;
    3602: romdata_int <= 'hb0d;
    3603: romdata_int <= 'h42d; // Line Descriptor
    3604: romdata_int <= 'h4200;
    3605: romdata_int <= 'h30c2;
    3606: romdata_int <= 'h1558;
    3607: romdata_int <= 'h42d; // Line Descriptor
    3608: romdata_int <= 'h4400;
    3609: romdata_int <= 'h48a4;
    3610: romdata_int <= 'h3354;
    3611: romdata_int <= 'h42d; // Line Descriptor
    3612: romdata_int <= 'h4600;
    3613: romdata_int <= 'h3a40;
    3614: romdata_int <= 'h3159;
    3615: romdata_int <= 'h42d; // Line Descriptor
    3616: romdata_int <= 'h4800;
    3617: romdata_int <= 'h3242;
    3618: romdata_int <= 'h2cb7;
    3619: romdata_int <= 'h42d; // Line Descriptor
    3620: romdata_int <= 'h4a00;
    3621: romdata_int <= 'h2d1;
    3622: romdata_int <= 'h2a6a;
    3623: romdata_int <= 'h42d; // Line Descriptor
    3624: romdata_int <= 'h4c00;
    3625: romdata_int <= 'h52f6;
    3626: romdata_int <= 'h4e6b;
    3627: romdata_int <= 'h42d; // Line Descriptor
    3628: romdata_int <= 'h4e00;
    3629: romdata_int <= 'h2c3e;
    3630: romdata_int <= 'h20bd;
    3631: romdata_int <= 'h42d; // Line Descriptor
    3632: romdata_int <= 'h5000;
    3633: romdata_int <= 'h20bc;
    3634: romdata_int <= 'h547;
    3635: romdata_int <= 'h42d; // Line Descriptor
    3636: romdata_int <= 'h5200;
    3637: romdata_int <= 'h46ad;
    3638: romdata_int <= 'h1f55;
    3639: romdata_int <= 'h42d; // Line Descriptor
    3640: romdata_int <= 'h5400;
    3641: romdata_int <= 'h121a;
    3642: romdata_int <= 'h26b0;
    3643: romdata_int <= 'h42d; // Line Descriptor
    3644: romdata_int <= 'h5600;
    3645: romdata_int <= 'h2234;
    3646: romdata_int <= 'h4cc0;
    3647: romdata_int <= 'h42d; // Line Descriptor
    3648: romdata_int <= 'h5800;
    3649: romdata_int <= 'h10ab;
    3650: romdata_int <= 'hc8a;
    3651: romdata_int <= 'h42d; // Line Descriptor
    3652: romdata_int <= 'h0;
    3653: romdata_int <= 'h184d;
    3654: romdata_int <= 'h49d;
    3655: romdata_int <= 'h42d; // Line Descriptor
    3656: romdata_int <= 'h200;
    3657: romdata_int <= 'h2057;
    3658: romdata_int <= 'h3d33;
    3659: romdata_int <= 'h42d; // Line Descriptor
    3660: romdata_int <= 'h400;
    3661: romdata_int <= 'h32aa;
    3662: romdata_int <= 'h3b1e;
    3663: romdata_int <= 'h42d; // Line Descriptor
    3664: romdata_int <= 'h600;
    3665: romdata_int <= 'h5826;
    3666: romdata_int <= 'h54b5;
    3667: romdata_int <= 'h42d; // Line Descriptor
    3668: romdata_int <= 'h800;
    3669: romdata_int <= 'had;
    3670: romdata_int <= 'ha1f;
    3671: romdata_int <= 'h42d; // Line Descriptor
    3672: romdata_int <= 'ha00;
    3673: romdata_int <= 'h42cc;
    3674: romdata_int <= 'h5282;
    3675: romdata_int <= 'h42d; // Line Descriptor
    3676: romdata_int <= 'hc00;
    3677: romdata_int <= 'h2637;
    3678: romdata_int <= 'h10ab;
    3679: romdata_int <= 'h42d; // Line Descriptor
    3680: romdata_int <= 'he00;
    3681: romdata_int <= 'h1639;
    3682: romdata_int <= 'h36af;
    3683: romdata_int <= 'h42d; // Line Descriptor
    3684: romdata_int <= 'h1000;
    3685: romdata_int <= 'hc6b;
    3686: romdata_int <= 'h2d5c;
    3687: romdata_int <= 'h42d; // Line Descriptor
    3688: romdata_int <= 'h1200;
    3689: romdata_int <= 'h3ee7;
    3690: romdata_int <= 'h1509;
    3691: romdata_int <= 'h42d; // Line Descriptor
    3692: romdata_int <= 'h1400;
    3693: romdata_int <= 'h1428;
    3694: romdata_int <= 'h814;
    3695: romdata_int <= 'h42d; // Line Descriptor
    3696: romdata_int <= 'h1600;
    3697: romdata_int <= 'h4afb;
    3698: romdata_int <= 'h4ecd;
    3699: romdata_int <= 'h42d; // Line Descriptor
    3700: romdata_int <= 'h1800;
    3701: romdata_int <= 'h22fb;
    3702: romdata_int <= 'h1e4f;
    3703: romdata_int <= 'h42d; // Line Descriptor
    3704: romdata_int <= 'h1a00;
    3705: romdata_int <= 'h2b4b;
    3706: romdata_int <= 'h503a;
    3707: romdata_int <= 'h42d; // Line Descriptor
    3708: romdata_int <= 'h1c00;
    3709: romdata_int <= 'h3aaa;
    3710: romdata_int <= 'h18ae;
    3711: romdata_int <= 'h42d; // Line Descriptor
    3712: romdata_int <= 'h1e00;
    3713: romdata_int <= 'h1c87;
    3714: romdata_int <= 'h4522;
    3715: romdata_int <= 'h42d; // Line Descriptor
    3716: romdata_int <= 'h2000;
    3717: romdata_int <= 'h2e57;
    3718: romdata_int <= 'hc3d;
    3719: romdata_int <= 'h42d; // Line Descriptor
    3720: romdata_int <= 'h2200;
    3721: romdata_int <= 'h8bd;
    3722: romdata_int <= 'h1a67;
    3723: romdata_int <= 'h42d; // Line Descriptor
    3724: romdata_int <= 'h2400;
    3725: romdata_int <= 'h130f;
    3726: romdata_int <= 'hec6;
    3727: romdata_int <= 'h42d; // Line Descriptor
    3728: romdata_int <= 'h2600;
    3729: romdata_int <= 'h447f;
    3730: romdata_int <= 'h2f14;
    3731: romdata_int <= 'h42d; // Line Descriptor
    3732: romdata_int <= 'h2800;
    3733: romdata_int <= 'h1b18;
    3734: romdata_int <= 'h2a62;
    3735: romdata_int <= 'h42d; // Line Descriptor
    3736: romdata_int <= 'h2a00;
    3737: romdata_int <= 'h4e1d;
    3738: romdata_int <= 'h1259;
    3739: romdata_int <= 'h42d; // Line Descriptor
    3740: romdata_int <= 'h2c00;
    3741: romdata_int <= 'h38bc;
    3742: romdata_int <= 'h4733;
    3743: romdata_int <= 'h42d; // Line Descriptor
    3744: romdata_int <= 'h2e00;
    3745: romdata_int <= 'h2826;
    3746: romdata_int <= 'h34b;
    3747: romdata_int <= 'h42d; // Line Descriptor
    3748: romdata_int <= 'h3000;
    3749: romdata_int <= 'h54c;
    3750: romdata_int <= 'h209e;
    3751: romdata_int <= 'h42d; // Line Descriptor
    3752: romdata_int <= 'h3200;
    3753: romdata_int <= 'h574c;
    3754: romdata_int <= 'h56c4;
    3755: romdata_int <= 'h42d; // Line Descriptor
    3756: romdata_int <= 'h3400;
    3757: romdata_int <= 'h1092;
    3758: romdata_int <= 'h1cbe;
    3759: romdata_int <= 'h42d; // Line Descriptor
    3760: romdata_int <= 'h3600;
    3761: romdata_int <= 'h546d;
    3762: romdata_int <= 'h4808;
    3763: romdata_int <= 'h42d; // Line Descriptor
    3764: romdata_int <= 'h3800;
    3765: romdata_int <= 'h3606;
    3766: romdata_int <= 'h331c;
    3767: romdata_int <= 'h42d; // Line Descriptor
    3768: romdata_int <= 'h3a00;
    3769: romdata_int <= 'h2534;
    3770: romdata_int <= 'h4094;
    3771: romdata_int <= 'h42d; // Line Descriptor
    3772: romdata_int <= 'h3c00;
    3773: romdata_int <= 'h2d07;
    3774: romdata_int <= 'h34f8;
    3775: romdata_int <= 'h42d; // Line Descriptor
    3776: romdata_int <= 'h3e00;
    3777: romdata_int <= 'h513f;
    3778: romdata_int <= 'h24ff;
    3779: romdata_int <= 'h42d; // Line Descriptor
    3780: romdata_int <= 'h4000;
    3781: romdata_int <= 'h4766;
    3782: romdata_int <= 'h1710;
    3783: romdata_int <= 'h42d; // Line Descriptor
    3784: romdata_int <= 'h4200;
    3785: romdata_int <= 'hf2b;
    3786: romdata_int <= 'h6a5;
    3787: romdata_int <= 'h42d; // Line Descriptor
    3788: romdata_int <= 'h4400;
    3789: romdata_int <= 'h4942;
    3790: romdata_int <= 'h3123;
    3791: romdata_int <= 'h42d; // Line Descriptor
    3792: romdata_int <= 'h4600;
    3793: romdata_int <= 'h1e38;
    3794: romdata_int <= 'h4cf9;
    3795: romdata_int <= 'h42d; // Line Descriptor
    3796: romdata_int <= 'h4800;
    3797: romdata_int <= 'h3c8f;
    3798: romdata_int <= 'h11a;
    3799: romdata_int <= 'h42d; // Line Descriptor
    3800: romdata_int <= 'h4a00;
    3801: romdata_int <= 'h4098;
    3802: romdata_int <= 'h26cf;
    3803: romdata_int <= 'h42d; // Line Descriptor
    3804: romdata_int <= 'h4c00;
    3805: romdata_int <= 'h3555;
    3806: romdata_int <= 'h3937;
    3807: romdata_int <= 'h42d; // Line Descriptor
    3808: romdata_int <= 'h4e00;
    3809: romdata_int <= 'h2b4;
    3810: romdata_int <= 'h22e2;
    3811: romdata_int <= 'h42d; // Line Descriptor
    3812: romdata_int <= 'h5000;
    3813: romdata_int <= 'h4d09;
    3814: romdata_int <= 'h426b;
    3815: romdata_int <= 'h42d; // Line Descriptor
    3816: romdata_int <= 'h5200;
    3817: romdata_int <= 'hb50;
    3818: romdata_int <= 'h5887;
    3819: romdata_int <= 'h42d; // Line Descriptor
    3820: romdata_int <= 'h5400;
    3821: romdata_int <= 'h52b2;
    3822: romdata_int <= 'h2941;
    3823: romdata_int <= 'h42d; // Line Descriptor
    3824: romdata_int <= 'h5600;
    3825: romdata_int <= 'h30f7;
    3826: romdata_int <= 'h4a72;
    3827: romdata_int <= 'h52d; // Line Descriptor
    3828: romdata_int <= 'h5800;
    3829: romdata_int <= 'h640;
    3830: romdata_int <= 'h3f42;
    3831: romdata_int <= 'h1424; // Line Descriptor
    3832: romdata_int <= 'h0;
    3833: romdata_int <= 'ha04;
    3834: romdata_int <= 'h2137;
    3835: romdata_int <= 'h3e9a;
    3836: romdata_int <= 'h30b0;
    3837: romdata_int <= 'h3f5c;
    3838: romdata_int <= 'h10e1;
    3839: romdata_int <= 'h12ec;
    3840: romdata_int <= 'h180b;
    3841: romdata_int <= 'h2516;
    3842: romdata_int <= 'h1964;
    3843: romdata_int <= 'h1424; // Line Descriptor
    3844: romdata_int <= 'h200;
    3845: romdata_int <= 'h2291;
    3846: romdata_int <= 'h2c0d;
    3847: romdata_int <= 'h2b28;
    3848: romdata_int <= 'h3c8a;
    3849: romdata_int <= 'h226b;
    3850: romdata_int <= 'h3467;
    3851: romdata_int <= 'h4055;
    3852: romdata_int <= 'h2261;
    3853: romdata_int <= 'h46d5;
    3854: romdata_int <= 'h131e;
    3855: romdata_int <= 'h1424; // Line Descriptor
    3856: romdata_int <= 'h400;
    3857: romdata_int <= 'h3cf2;
    3858: romdata_int <= 'h129a;
    3859: romdata_int <= 'h184e;
    3860: romdata_int <= 'h3ac4;
    3861: romdata_int <= 'h2950;
    3862: romdata_int <= 'h1323;
    3863: romdata_int <= 'h300f;
    3864: romdata_int <= 'h26d8;
    3865: romdata_int <= 'h2852;
    3866: romdata_int <= 'h423b;
    3867: romdata_int <= 'h1424; // Line Descriptor
    3868: romdata_int <= 'h600;
    3869: romdata_int <= 'h464a;
    3870: romdata_int <= 'h2877;
    3871: romdata_int <= 'h44e7;
    3872: romdata_int <= 'h3813;
    3873: romdata_int <= 'h424e;
    3874: romdata_int <= 'h145a;
    3875: romdata_int <= 'h1e83;
    3876: romdata_int <= 'h3318;
    3877: romdata_int <= 'h1a0e;
    3878: romdata_int <= 'h38d0;
    3879: romdata_int <= 'h1424; // Line Descriptor
    3880: romdata_int <= 'h800;
    3881: romdata_int <= 'hf4f;
    3882: romdata_int <= 'h2625;
    3883: romdata_int <= 'h94d;
    3884: romdata_int <= 'h2f52;
    3885: romdata_int <= 'h4738;
    3886: romdata_int <= 'h1a8f;
    3887: romdata_int <= 'h420e;
    3888: romdata_int <= 'h14ab;
    3889: romdata_int <= 'h4475;
    3890: romdata_int <= 'h2e41;
    3891: romdata_int <= 'h1424; // Line Descriptor
    3892: romdata_int <= 'ha00;
    3893: romdata_int <= 'h30bd;
    3894: romdata_int <= 'h1ec5;
    3895: romdata_int <= 'h63b;
    3896: romdata_int <= 'h2067;
    3897: romdata_int <= 'h269f;
    3898: romdata_int <= 'h3132;
    3899: romdata_int <= 'h392a;
    3900: romdata_int <= 'ha71;
    3901: romdata_int <= 'h61c;
    3902: romdata_int <= 'h45f;
    3903: romdata_int <= 'h1424; // Line Descriptor
    3904: romdata_int <= 'hc00;
    3905: romdata_int <= 'h3738;
    3906: romdata_int <= 'h3821;
    3907: romdata_int <= 'h2d08;
    3908: romdata_int <= 'h3428;
    3909: romdata_int <= 'h212c;
    3910: romdata_int <= 'h81a;
    3911: romdata_int <= 'h68;
    3912: romdata_int <= 'he4e;
    3913: romdata_int <= 'h2d3f;
    3914: romdata_int <= 'h2341;
    3915: romdata_int <= 'h1424; // Line Descriptor
    3916: romdata_int <= 'he00;
    3917: romdata_int <= 'h1a7e;
    3918: romdata_int <= 'h2f3f;
    3919: romdata_int <= 'h41f;
    3920: romdata_int <= 'h1c23;
    3921: romdata_int <= 'h1f46;
    3922: romdata_int <= 'h2e90;
    3923: romdata_int <= 'hcda;
    3924: romdata_int <= 'h2f63;
    3925: romdata_int <= 'h1e70;
    3926: romdata_int <= 'h8b4;
    3927: romdata_int <= 'h1424; // Line Descriptor
    3928: romdata_int <= 'h1000;
    3929: romdata_int <= 'hcea;
    3930: romdata_int <= 'h1672;
    3931: romdata_int <= 'h1106;
    3932: romdata_int <= 'h220b;
    3933: romdata_int <= 'h367b;
    3934: romdata_int <= 'h3c3e;
    3935: romdata_int <= 'h3edb;
    3936: romdata_int <= 'h2558;
    3937: romdata_int <= 'h16ee;
    3938: romdata_int <= 'h40c3;
    3939: romdata_int <= 'h1424; // Line Descriptor
    3940: romdata_int <= 'h1200;
    3941: romdata_int <= 'h426b;
    3942: romdata_int <= 'h24fd;
    3943: romdata_int <= 'h1a9d;
    3944: romdata_int <= 'ha7d;
    3945: romdata_int <= 'h641;
    3946: romdata_int <= 'h207;
    3947: romdata_int <= 'h3682;
    3948: romdata_int <= 'h4467;
    3949: romdata_int <= 'h3473;
    3950: romdata_int <= 'h102b;
    3951: romdata_int <= 'h1424; // Line Descriptor
    3952: romdata_int <= 'h1400;
    3953: romdata_int <= 'h182f;
    3954: romdata_int <= 'h10f8;
    3955: romdata_int <= 'hebc;
    3956: romdata_int <= 'h46ef;
    3957: romdata_int <= 'hee3;
    3958: romdata_int <= 'h44dc;
    3959: romdata_int <= 'h34e4;
    3960: romdata_int <= 'h4da;
    3961: romdata_int <= 'h36f6;
    3962: romdata_int <= 'h2f2;
    3963: romdata_int <= 'h1424; // Line Descriptor
    3964: romdata_int <= 'h1600;
    3965: romdata_int <= 'h2145;
    3966: romdata_int <= 'h3078;
    3967: romdata_int <= 'h1efc;
    3968: romdata_int <= 'h4138;
    3969: romdata_int <= 'hc3f;
    3970: romdata_int <= 'h18f5;
    3971: romdata_int <= 'h6fe;
    3972: romdata_int <= 'h1d4b;
    3973: romdata_int <= 'hca8;
    3974: romdata_int <= 'h2697;
    3975: romdata_int <= 'h1424; // Line Descriptor
    3976: romdata_int <= 'h1800;
    3977: romdata_int <= 'h1ecb;
    3978: romdata_int <= 'h146e;
    3979: romdata_int <= 'h431e;
    3980: romdata_int <= 'h143c;
    3981: romdata_int <= 'h24e5;
    3982: romdata_int <= 'h46b;
    3983: romdata_int <= 'h4639;
    3984: romdata_int <= 'h1766;
    3985: romdata_int <= 'h3b07;
    3986: romdata_int <= 'h145;
    3987: romdata_int <= 'h1424; // Line Descriptor
    3988: romdata_int <= 'h1a00;
    3989: romdata_int <= 'h347a;
    3990: romdata_int <= 'h3628;
    3991: romdata_int <= 'hc45;
    3992: romdata_int <= 'h12a2;
    3993: romdata_int <= 'h3216;
    3994: romdata_int <= 'hb3e;
    3995: romdata_int <= 'h3a0e;
    3996: romdata_int <= 'h2b37;
    3997: romdata_int <= 'h154c;
    3998: romdata_int <= 'h3e91;
    3999: romdata_int <= 'h1424; // Line Descriptor
    4000: romdata_int <= 'h1c00;
    4001: romdata_int <= 'h3a2a;
    4002: romdata_int <= 'h327d;
    4003: romdata_int <= 'h28dd;
    4004: romdata_int <= 'h260;
    4005: romdata_int <= 'h4108;
    4006: romdata_int <= 'h2ad6;
    4007: romdata_int <= 'h1069;
    4008: romdata_int <= 'h3c52;
    4009: romdata_int <= 'heaf;
    4010: romdata_int <= 'h2aa6;
    4011: romdata_int <= 'h1424; // Line Descriptor
    4012: romdata_int <= 'h1e00;
    4013: romdata_int <= 'h13f;
    4014: romdata_int <= 'h64c;
    4015: romdata_int <= 'h366f;
    4016: romdata_int <= 'h1750;
    4017: romdata_int <= 'hb5;
    4018: romdata_int <= 'h160f;
    4019: romdata_int <= 'h2047;
    4020: romdata_int <= 'h8b8;
    4021: romdata_int <= 'h1ce2;
    4022: romdata_int <= 'h3111;
    4023: romdata_int <= 'h1424; // Line Descriptor
    4024: romdata_int <= 'h2000;
    4025: romdata_int <= 'h2ca8;
    4026: romdata_int <= 'h4230;
    4027: romdata_int <= 'h2680;
    4028: romdata_int <= 'h24b5;
    4029: romdata_int <= 'h3adb;
    4030: romdata_int <= 'h2c67;
    4031: romdata_int <= 'h2d49;
    4032: romdata_int <= 'h1a32;
    4033: romdata_int <= 'h3d55;
    4034: romdata_int <= 'hae5;
    4035: romdata_int <= 'h1424; // Line Descriptor
    4036: romdata_int <= 'h2200;
    4037: romdata_int <= 'h2b59;
    4038: romdata_int <= 'h2298;
    4039: romdata_int <= 'hf3;
    4040: romdata_int <= 'h32d9;
    4041: romdata_int <= 'h38d4;
    4042: romdata_int <= 'h1c3a;
    4043: romdata_int <= 'h33b;
    4044: romdata_int <= 'h2851;
    4045: romdata_int <= 'h20ba;
    4046: romdata_int <= 'h334c;
    4047: romdata_int <= 'h424; // Line Descriptor
    4048: romdata_int <= 'h2400;
    4049: romdata_int <= 'h71a;
    4050: romdata_int <= 'h4474;
    4051: romdata_int <= 'h424; // Line Descriptor
    4052: romdata_int <= 'h2600;
    4053: romdata_int <= 'h41c;
    4054: romdata_int <= 'hf23;
    4055: romdata_int <= 'h424; // Line Descriptor
    4056: romdata_int <= 'h2800;
    4057: romdata_int <= 'h10f7;
    4058: romdata_int <= 'h351c;
    4059: romdata_int <= 'h424; // Line Descriptor
    4060: romdata_int <= 'h2a00;
    4061: romdata_int <= 'h271c;
    4062: romdata_int <= 'h555;
    4063: romdata_int <= 'h424; // Line Descriptor
    4064: romdata_int <= 'h2c00;
    4065: romdata_int <= 'h1cc4;
    4066: romdata_int <= 'ha7a;
    4067: romdata_int <= 'h424; // Line Descriptor
    4068: romdata_int <= 'h2e00;
    4069: romdata_int <= 'h3f54;
    4070: romdata_int <= 'h466b;
    4071: romdata_int <= 'h424; // Line Descriptor
    4072: romdata_int <= 'h3000;
    4073: romdata_int <= 'h394c;
    4074: romdata_int <= 'h40bd;
    4075: romdata_int <= 'h424; // Line Descriptor
    4076: romdata_int <= 'h3200;
    4077: romdata_int <= 'h1508;
    4078: romdata_int <= 'h79;
    4079: romdata_int <= 'h424; // Line Descriptor
    4080: romdata_int <= 'h3400;
    4081: romdata_int <= 'h12c6;
    4082: romdata_int <= 'h2b1d;
    4083: romdata_int <= 'h424; // Line Descriptor
    4084: romdata_int <= 'h3600;
    4085: romdata_int <= 'h34a;
    4086: romdata_int <= 'hc46;
    4087: romdata_int <= 'h424; // Line Descriptor
    4088: romdata_int <= 'h3800;
    4089: romdata_int <= 'h3236;
    4090: romdata_int <= 'h3b3e;
    4091: romdata_int <= 'h424; // Line Descriptor
    4092: romdata_int <= 'h3a00;
    4093: romdata_int <= 'h2854;
    4094: romdata_int <= 'h1b2f;
    4095: romdata_int <= 'h424; // Line Descriptor
    4096: romdata_int <= 'h3c00;
    4097: romdata_int <= 'h83e;
    4098: romdata_int <= 'h18f2;
    4099: romdata_int <= 'h424; // Line Descriptor
    4100: romdata_int <= 'h3e00;
    4101: romdata_int <= 'h40fc;
    4102: romdata_int <= 'h8b0;
    4103: romdata_int <= 'h424; // Line Descriptor
    4104: romdata_int <= 'h4000;
    4105: romdata_int <= 'h44cb;
    4106: romdata_int <= 'h1cee;
    4107: romdata_int <= 'h424; // Line Descriptor
    4108: romdata_int <= 'h4200;
    4109: romdata_int <= 'h1744;
    4110: romdata_int <= 'h321;
    4111: romdata_int <= 'h424; // Line Descriptor
    4112: romdata_int <= 'h4400;
    4113: romdata_int <= 'h2eb3;
    4114: romdata_int <= 'h3f62;
    4115: romdata_int <= 'h424; // Line Descriptor
    4116: romdata_int <= 'h4600;
    4117: romdata_int <= 'h2458;
    4118: romdata_int <= 'h3d52;
    4119: romdata_int <= 'h424; // Line Descriptor
    4120: romdata_int <= 'h0;
    4121: romdata_int <= 'h130b;
    4122: romdata_int <= 'h433d;
    4123: romdata_int <= 'h424; // Line Descriptor
    4124: romdata_int <= 'h200;
    4125: romdata_int <= 'h44cf;
    4126: romdata_int <= 'h3e9b;
    4127: romdata_int <= 'h424; // Line Descriptor
    4128: romdata_int <= 'h400;
    4129: romdata_int <= 'h4677;
    4130: romdata_int <= 'h2687;
    4131: romdata_int <= 'h424; // Line Descriptor
    4132: romdata_int <= 'h600;
    4133: romdata_int <= 'h3d;
    4134: romdata_int <= 'h2809;
    4135: romdata_int <= 'h424; // Line Descriptor
    4136: romdata_int <= 'h800;
    4137: romdata_int <= 'h6d1;
    4138: romdata_int <= 'h34b8;
    4139: romdata_int <= 'h424; // Line Descriptor
    4140: romdata_int <= 'ha00;
    4141: romdata_int <= 'h329;
    4142: romdata_int <= 'h3843;
    4143: romdata_int <= 'h424; // Line Descriptor
    4144: romdata_int <= 'hc00;
    4145: romdata_int <= 'h2ebb;
    4146: romdata_int <= 'hc4b;
    4147: romdata_int <= 'h424; // Line Descriptor
    4148: romdata_int <= 'he00;
    4149: romdata_int <= 'h408e;
    4150: romdata_int <= 'h2ca6;
    4151: romdata_int <= 'h424; // Line Descriptor
    4152: romdata_int <= 'h1000;
    4153: romdata_int <= 'h3732;
    4154: romdata_int <= 'hadf;
    4155: romdata_int <= 'h424; // Line Descriptor
    4156: romdata_int <= 'h1200;
    4157: romdata_int <= 'h2c86;
    4158: romdata_int <= 'he7b;
    4159: romdata_int <= 'h424; // Line Descriptor
    4160: romdata_int <= 'h1400;
    4161: romdata_int <= 'h2273;
    4162: romdata_int <= 'h1900;
    4163: romdata_int <= 'h424; // Line Descriptor
    4164: romdata_int <= 'h1600;
    4165: romdata_int <= 'h3d54;
    4166: romdata_int <= 'h14b6;
    4167: romdata_int <= 'h424; // Line Descriptor
    4168: romdata_int <= 'h1800;
    4169: romdata_int <= 'h54c;
    4170: romdata_int <= 'h40d2;
    4171: romdata_int <= 'h424; // Line Descriptor
    4172: romdata_int <= 'h1a00;
    4173: romdata_int <= 'h8ce;
    4174: romdata_int <= 'h48;
    4175: romdata_int <= 'h424; // Line Descriptor
    4176: romdata_int <= 'h1c00;
    4177: romdata_int <= 'h34f4;
    4178: romdata_int <= 'h310b;
    4179: romdata_int <= 'h424; // Line Descriptor
    4180: romdata_int <= 'h1e00;
    4181: romdata_int <= 'ha13;
    4182: romdata_int <= 'h3c96;
    4183: romdata_int <= 'h424; // Line Descriptor
    4184: romdata_int <= 'h2000;
    4185: romdata_int <= 'h2819;
    4186: romdata_int <= 'h1024;
    4187: romdata_int <= 'h424; // Line Descriptor
    4188: romdata_int <= 'h2200;
    4189: romdata_int <= 'h3a22;
    4190: romdata_int <= 'h254b;
    4191: romdata_int <= 'h424; // Line Descriptor
    4192: romdata_int <= 'h2400;
    4193: romdata_int <= 'h2709;
    4194: romdata_int <= 'h8a7;
    4195: romdata_int <= 'h424; // Line Descriptor
    4196: romdata_int <= 'h2600;
    4197: romdata_int <= 'h3008;
    4198: romdata_int <= 'h3ad2;
    4199: romdata_int <= 'h424; // Line Descriptor
    4200: romdata_int <= 'h2800;
    4201: romdata_int <= 'h167b;
    4202: romdata_int <= 'h2a74;
    4203: romdata_int <= 'h424; // Line Descriptor
    4204: romdata_int <= 'h2a00;
    4205: romdata_int <= 'hc6f;
    4206: romdata_int <= 'h1f09;
    4207: romdata_int <= 'h424; // Line Descriptor
    4208: romdata_int <= 'h2c00;
    4209: romdata_int <= 'h3953;
    4210: romdata_int <= 'h6d8;
    4211: romdata_int <= 'h424; // Line Descriptor
    4212: romdata_int <= 'h2e00;
    4213: romdata_int <= 'h2429;
    4214: romdata_int <= 'h44f3;
    4215: romdata_int <= 'h424; // Line Descriptor
    4216: romdata_int <= 'h3000;
    4217: romdata_int <= 'h2b2a;
    4218: romdata_int <= 'h126e;
    4219: romdata_int <= 'h424; // Line Descriptor
    4220: romdata_int <= 'h3200;
    4221: romdata_int <= 'h1879;
    4222: romdata_int <= 'h2e60;
    4223: romdata_int <= 'h424; // Line Descriptor
    4224: romdata_int <= 'h3400;
    4225: romdata_int <= 'h20af;
    4226: romdata_int <= 'h1c94;
    4227: romdata_int <= 'h424; // Line Descriptor
    4228: romdata_int <= 'h3600;
    4229: romdata_int <= 'he44;
    4230: romdata_int <= 'h261;
    4231: romdata_int <= 'h424; // Line Descriptor
    4232: romdata_int <= 'h3800;
    4233: romdata_int <= 'h3351;
    4234: romdata_int <= 'h32cd;
    4235: romdata_int <= 'h424; // Line Descriptor
    4236: romdata_int <= 'h3a00;
    4237: romdata_int <= 'h14b7;
    4238: romdata_int <= 'h173f;
    4239: romdata_int <= 'h424; // Line Descriptor
    4240: romdata_int <= 'h3c00;
    4241: romdata_int <= 'h4347;
    4242: romdata_int <= 'h367b;
    4243: romdata_int <= 'h424; // Line Descriptor
    4244: romdata_int <= 'h3e00;
    4245: romdata_int <= 'h1b0b;
    4246: romdata_int <= 'h43a;
    4247: romdata_int <= 'h424; // Line Descriptor
    4248: romdata_int <= 'h4000;
    4249: romdata_int <= 'h1e83;
    4250: romdata_int <= 'h2240;
    4251: romdata_int <= 'h424; // Line Descriptor
    4252: romdata_int <= 'h4200;
    4253: romdata_int <= 'h1c63;
    4254: romdata_int <= 'h2048;
    4255: romdata_int <= 'h424; // Line Descriptor
    4256: romdata_int <= 'h4400;
    4257: romdata_int <= 'h10ec;
    4258: romdata_int <= 'h1a33;
    4259: romdata_int <= 'h424; // Line Descriptor
    4260: romdata_int <= 'h4600;
    4261: romdata_int <= 'h3e6f;
    4262: romdata_int <= 'h461f;
    4263: romdata_int <= 'h424; // Line Descriptor
    4264: romdata_int <= 'h0;
    4265: romdata_int <= 'h3e9c;
    4266: romdata_int <= 'h689;
    4267: romdata_int <= 'h424; // Line Descriptor
    4268: romdata_int <= 'h200;
    4269: romdata_int <= 'he75;
    4270: romdata_int <= 'h4433;
    4271: romdata_int <= 'h424; // Line Descriptor
    4272: romdata_int <= 'h400;
    4273: romdata_int <= 'h3130;
    4274: romdata_int <= 'h34df;
    4275: romdata_int <= 'h424; // Line Descriptor
    4276: romdata_int <= 'h600;
    4277: romdata_int <= 'h2cc1;
    4278: romdata_int <= 'h1697;
    4279: romdata_int <= 'h424; // Line Descriptor
    4280: romdata_int <= 'h800;
    4281: romdata_int <= 'h1a59;
    4282: romdata_int <= 'h2c9c;
    4283: romdata_int <= 'h424; // Line Descriptor
    4284: romdata_int <= 'ha00;
    4285: romdata_int <= 'h10f9;
    4286: romdata_int <= 'h2a12;
    4287: romdata_int <= 'h424; // Line Descriptor
    4288: romdata_int <= 'hc00;
    4289: romdata_int <= 'h49c;
    4290: romdata_int <= 'h215a;
    4291: romdata_int <= 'h424; // Line Descriptor
    4292: romdata_int <= 'he00;
    4293: romdata_int <= 'h2228;
    4294: romdata_int <= 'h2823;
    4295: romdata_int <= 'h424; // Line Descriptor
    4296: romdata_int <= 'h1000;
    4297: romdata_int <= 'h18f6;
    4298: romdata_int <= 'h3e6b;
    4299: romdata_int <= 'h424; // Line Descriptor
    4300: romdata_int <= 'h1200;
    4301: romdata_int <= 'h14f6;
    4302: romdata_int <= 'h22;
    4303: romdata_int <= 'h424; // Line Descriptor
    4304: romdata_int <= 'h1400;
    4305: romdata_int <= 'h26e8;
    4306: romdata_int <= 'h40a5;
    4307: romdata_int <= 'h424; // Line Descriptor
    4308: romdata_int <= 'h1600;
    4309: romdata_int <= 'h1c07;
    4310: romdata_int <= 'h1a7a;
    4311: romdata_int <= 'h424; // Line Descriptor
    4312: romdata_int <= 'h1800;
    4313: romdata_int <= 'h4466;
    4314: romdata_int <= 'h85a;
    4315: romdata_int <= 'h424; // Line Descriptor
    4316: romdata_int <= 'h1a00;
    4317: romdata_int <= 'h36a7;
    4318: romdata_int <= 'h18a2;
    4319: romdata_int <= 'h424; // Line Descriptor
    4320: romdata_int <= 'h1c00;
    4321: romdata_int <= 'hc8;
    4322: romdata_int <= 'he5b;
    4323: romdata_int <= 'h424; // Line Descriptor
    4324: romdata_int <= 'h1e00;
    4325: romdata_int <= 'h3429;
    4326: romdata_int <= 'h1d39;
    4327: romdata_int <= 'h424; // Line Descriptor
    4328: romdata_int <= 'h2000;
    4329: romdata_int <= 'hd56;
    4330: romdata_int <= 'hc3d;
    4331: romdata_int <= 'h424; // Line Descriptor
    4332: romdata_int <= 'h2200;
    4333: romdata_int <= 'h2e7d;
    4334: romdata_int <= 'h3a1a;
    4335: romdata_int <= 'h424; // Line Descriptor
    4336: romdata_int <= 'h2400;
    4337: romdata_int <= 'h170a;
    4338: romdata_int <= 'h36c2;
    4339: romdata_int <= 'h424; // Line Descriptor
    4340: romdata_int <= 'h2600;
    4341: romdata_int <= 'h4046;
    4342: romdata_int <= 'h4638;
    4343: romdata_int <= 'h424; // Line Descriptor
    4344: romdata_int <= 'h2800;
    4345: romdata_int <= 'h2b4e;
    4346: romdata_int <= 'h151e;
    4347: romdata_int <= 'h424; // Line Descriptor
    4348: romdata_int <= 'h2a00;
    4349: romdata_int <= 'h2533;
    4350: romdata_int <= 'h388d;
    4351: romdata_int <= 'h424; // Line Descriptor
    4352: romdata_int <= 'h2c00;
    4353: romdata_int <= 'h6b8;
    4354: romdata_int <= 'h3cbf;
    4355: romdata_int <= 'h424; // Line Descriptor
    4356: romdata_int <= 'h2e00;
    4357: romdata_int <= 'h3312;
    4358: romdata_int <= 'h423a;
    4359: romdata_int <= 'h424; // Line Descriptor
    4360: romdata_int <= 'h3000;
    4361: romdata_int <= 'h217;
    4362: romdata_int <= 'h230d;
    4363: romdata_int <= 'h424; // Line Descriptor
    4364: romdata_int <= 'h3200;
    4365: romdata_int <= 'ha3d;
    4366: romdata_int <= 'h2632;
    4367: romdata_int <= 'h424; // Line Descriptor
    4368: romdata_int <= 'h3400;
    4369: romdata_int <= 'h3ab9;
    4370: romdata_int <= 'h367;
    4371: romdata_int <= 'h424; // Line Descriptor
    4372: romdata_int <= 'h3600;
    4373: romdata_int <= 'h1e3b;
    4374: romdata_int <= 'h12f3;
    4375: romdata_int <= 'h424; // Line Descriptor
    4376: romdata_int <= 'h3800;
    4377: romdata_int <= 'h214d;
    4378: romdata_int <= 'h10a5;
    4379: romdata_int <= 'h424; // Line Descriptor
    4380: romdata_int <= 'h3a00;
    4381: romdata_int <= 'h38f1;
    4382: romdata_int <= 'h2e58;
    4383: romdata_int <= 'h424; // Line Descriptor
    4384: romdata_int <= 'h3c00;
    4385: romdata_int <= 'h46e2;
    4386: romdata_int <= 'h332f;
    4387: romdata_int <= 'h424; // Line Descriptor
    4388: romdata_int <= 'h3e00;
    4389: romdata_int <= 'h42ae;
    4390: romdata_int <= 'h30c5;
    4391: romdata_int <= 'h424; // Line Descriptor
    4392: romdata_int <= 'h4000;
    4393: romdata_int <= 'h811;
    4394: romdata_int <= 'h24c6;
    4395: romdata_int <= 'h424; // Line Descriptor
    4396: romdata_int <= 'h4200;
    4397: romdata_int <= 'h3c8e;
    4398: romdata_int <= 'hb0f;
    4399: romdata_int <= 'h424; // Line Descriptor
    4400: romdata_int <= 'h4400;
    4401: romdata_int <= 'h1320;
    4402: romdata_int <= 'h4e2;
    4403: romdata_int <= 'h424; // Line Descriptor
    4404: romdata_int <= 'h4600;
    4405: romdata_int <= 'h28d3;
    4406: romdata_int <= 'h1ea1;
    4407: romdata_int <= 'h424; // Line Descriptor
    4408: romdata_int <= 'h0;
    4409: romdata_int <= 'h1aca;
    4410: romdata_int <= 'h4711;
    4411: romdata_int <= 'h424; // Line Descriptor
    4412: romdata_int <= 'h200;
    4413: romdata_int <= 'h30d7;
    4414: romdata_int <= 'h3f2d;
    4415: romdata_int <= 'h424; // Line Descriptor
    4416: romdata_int <= 'h400;
    4417: romdata_int <= 'h3f56;
    4418: romdata_int <= 'h26fa;
    4419: romdata_int <= 'h424; // Line Descriptor
    4420: romdata_int <= 'h600;
    4421: romdata_int <= 'h2c7a;
    4422: romdata_int <= 'h1ee7;
    4423: romdata_int <= 'h424; // Line Descriptor
    4424: romdata_int <= 'h800;
    4425: romdata_int <= 'h1060;
    4426: romdata_int <= 'h3c11;
    4427: romdata_int <= 'h424; // Line Descriptor
    4428: romdata_int <= 'ha00;
    4429: romdata_int <= 'h18c1;
    4430: romdata_int <= 'h2e38;
    4431: romdata_int <= 'h424; // Line Descriptor
    4432: romdata_int <= 'hc00;
    4433: romdata_int <= 'h3c15;
    4434: romdata_int <= 'h4253;
    4435: romdata_int <= 'h424; // Line Descriptor
    4436: romdata_int <= 'he00;
    4437: romdata_int <= 'h3413;
    4438: romdata_int <= 'h4439;
    4439: romdata_int <= 'h424; // Line Descriptor
    4440: romdata_int <= 'h1000;
    4441: romdata_int <= 'hece;
    4442: romdata_int <= 'h2a9b;
    4443: romdata_int <= 'h424; // Line Descriptor
    4444: romdata_int <= 'h1200;
    4445: romdata_int <= 'h28e1;
    4446: romdata_int <= 'h3287;
    4447: romdata_int <= 'h424; // Line Descriptor
    4448: romdata_int <= 'h1400;
    4449: romdata_int <= 'h358;
    4450: romdata_int <= 'h54d;
    4451: romdata_int <= 'h424; // Line Descriptor
    4452: romdata_int <= 'h1600;
    4453: romdata_int <= 'h270e;
    4454: romdata_int <= 'h3516;
    4455: romdata_int <= 'h424; // Line Descriptor
    4456: romdata_int <= 'h1800;
    4457: romdata_int <= 'h380b;
    4458: romdata_int <= 'h151a;
    4459: romdata_int <= 'h424; // Line Descriptor
    4460: romdata_int <= 'h1a00;
    4461: romdata_int <= 'h1e25;
    4462: romdata_int <= 'h2d3;
    4463: romdata_int <= 'h424; // Line Descriptor
    4464: romdata_int <= 'h1c00;
    4465: romdata_int <= 'h1428;
    4466: romdata_int <= 'h803;
    4467: romdata_int <= 'h424; // Line Descriptor
    4468: romdata_int <= 'h1e00;
    4469: romdata_int <= 'h12dd;
    4470: romdata_int <= 'h24eb;
    4471: romdata_int <= 'h424; // Line Descriptor
    4472: romdata_int <= 'h2000;
    4473: romdata_int <= 'h22f8;
    4474: romdata_int <= 'h22cd;
    4475: romdata_int <= 'h424; // Line Descriptor
    4476: romdata_int <= 'h2200;
    4477: romdata_int <= 'h4b7;
    4478: romdata_int <= 'he7;
    4479: romdata_int <= 'h424; // Line Descriptor
    4480: romdata_int <= 'h2400;
    4481: romdata_int <= 'h44bd;
    4482: romdata_int <= 'h16fa;
    4483: romdata_int <= 'h424; // Line Descriptor
    4484: romdata_int <= 'h2600;
    4485: romdata_int <= 'h24ab;
    4486: romdata_int <= 'h1d05;
    4487: romdata_int <= 'h424; // Line Descriptor
    4488: romdata_int <= 'h2800;
    4489: romdata_int <= 'h607;
    4490: romdata_int <= 'ha03;
    4491: romdata_int <= 'h424; // Line Descriptor
    4492: romdata_int <= 'h2a00;
    4493: romdata_int <= 'haac;
    4494: romdata_int <= 'h6a2;
    4495: romdata_int <= 'h424; // Line Descriptor
    4496: romdata_int <= 'h2c00;
    4497: romdata_int <= 'h1d66;
    4498: romdata_int <= 'h386a;
    4499: romdata_int <= 'h424; // Line Descriptor
    4500: romdata_int <= 'h2e00;
    4501: romdata_int <= 'h2a79;
    4502: romdata_int <= 'h1a61;
    4503: romdata_int <= 'h424; // Line Descriptor
    4504: romdata_int <= 'h3000;
    4505: romdata_int <= 'hc98;
    4506: romdata_int <= 'h40f0;
    4507: romdata_int <= 'h424; // Line Descriptor
    4508: romdata_int <= 'h3200;
    4509: romdata_int <= 'h327b;
    4510: romdata_int <= 'h103b;
    4511: romdata_int <= 'h424; // Line Descriptor
    4512: romdata_int <= 'h3400;
    4513: romdata_int <= 'h90e;
    4514: romdata_int <= 'h1826;
    4515: romdata_int <= 'h424; // Line Descriptor
    4516: romdata_int <= 'h3600;
    4517: romdata_int <= 'h4750;
    4518: romdata_int <= 'hd40;
    4519: romdata_int <= 'h424; // Line Descriptor
    4520: romdata_int <= 'h3800;
    4521: romdata_int <= 'h1756;
    4522: romdata_int <= 'hf08;
    4523: romdata_int <= 'h424; // Line Descriptor
    4524: romdata_int <= 'h3a00;
    4525: romdata_int <= 'h2ee4;
    4526: romdata_int <= 'h3030;
    4527: romdata_int <= 'h424; // Line Descriptor
    4528: romdata_int <= 'h3c00;
    4529: romdata_int <= 'h3a0d;
    4530: romdata_int <= 'h2cfa;
    4531: romdata_int <= 'h424; // Line Descriptor
    4532: romdata_int <= 'h3e00;
    4533: romdata_int <= 'h102;
    4534: romdata_int <= 'h2855;
    4535: romdata_int <= 'h424; // Line Descriptor
    4536: romdata_int <= 'h4000;
    4537: romdata_int <= 'h4244;
    4538: romdata_int <= 'h36d0;
    4539: romdata_int <= 'h424; // Line Descriptor
    4540: romdata_int <= 'h4200;
    4541: romdata_int <= 'h404a;
    4542: romdata_int <= 'h2007;
    4543: romdata_int <= 'h424; // Line Descriptor
    4544: romdata_int <= 'h4400;
    4545: romdata_int <= 'h366f;
    4546: romdata_int <= 'h3b56;
    4547: romdata_int <= 'h524; // Line Descriptor
    4548: romdata_int <= 'h4600;
    4549: romdata_int <= 'h20c5;
    4550: romdata_int <= 'h129a;
    4551: romdata_int <= 'h181e; // Line Descriptor
    4552: romdata_int <= 'h0;
    4553: romdata_int <= 'h1891;
    4554: romdata_int <= 'h340d;
    4555: romdata_int <= 'h3b28;
    4556: romdata_int <= 'h208a;
    4557: romdata_int <= 'hc6b;
    4558: romdata_int <= 'h2c67;
    4559: romdata_int <= 'h1455;
    4560: romdata_int <= 'h461;
    4561: romdata_int <= 'h1ed5;
    4562: romdata_int <= 'h1b1e;
    4563: romdata_int <= 'h26a5;
    4564: romdata_int <= 'h6e0;
    4565: romdata_int <= 'h181e; // Line Descriptor
    4566: romdata_int <= 'h200;
    4567: romdata_int <= 'h2652;
    4568: romdata_int <= 'h203b;
    4569: romdata_int <= 'h112b;
    4570: romdata_int <= 'h1664;
    4571: romdata_int <= 'h2690;
    4572: romdata_int <= 'h1b36;
    4573: romdata_int <= 'hed5;
    4574: romdata_int <= 'h2262;
    4575: romdata_int <= 'h38f2;
    4576: romdata_int <= 'h30b6;
    4577: romdata_int <= 'h2c9;
    4578: romdata_int <= 'h2354;
    4579: romdata_int <= 'h181e; // Line Descriptor
    4580: romdata_int <= 'h400;
    4581: romdata_int <= 'hb53;
    4582: romdata_int <= 'h132c;
    4583: romdata_int <= 'h2749;
    4584: romdata_int <= 'h267;
    4585: romdata_int <= 'haa6;
    4586: romdata_int <= 'hef2;
    4587: romdata_int <= 'h1888;
    4588: romdata_int <= 'h3127;
    4589: romdata_int <= 'h2bd;
    4590: romdata_int <= 'h225c;
    4591: romdata_int <= 'h3a48;
    4592: romdata_int <= 'h2122;
    4593: romdata_int <= 'h181e; // Line Descriptor
    4594: romdata_int <= 'h600;
    4595: romdata_int <= 'h2d2d;
    4596: romdata_int <= 'h329f;
    4597: romdata_int <= 'h3082;
    4598: romdata_int <= 'h1470;
    4599: romdata_int <= 'h114f;
    4600: romdata_int <= 'h2425;
    4601: romdata_int <= 'hd4d;
    4602: romdata_int <= 'h3352;
    4603: romdata_int <= 'h138;
    4604: romdata_int <= 'he8f;
    4605: romdata_int <= 'h1c0e;
    4606: romdata_int <= 'h10ab;
    4607: romdata_int <= 'h181e; // Line Descriptor
    4608: romdata_int <= 'h800;
    4609: romdata_int <= 'h124f;
    4610: romdata_int <= 'h905;
    4611: romdata_int <= 'haa1;
    4612: romdata_int <= 'h224d;
    4613: romdata_int <= 'h748;
    4614: romdata_int <= 'h301a;
    4615: romdata_int <= 'h3a0a;
    4616: romdata_int <= 'h1b16;
    4617: romdata_int <= 'h36ee;
    4618: romdata_int <= 'h1466;
    4619: romdata_int <= 'h3832;
    4620: romdata_int <= 'h2af3;
    4621: romdata_int <= 'h181e; // Line Descriptor
    4622: romdata_int <= 'ha00;
    4623: romdata_int <= 'h1e72;
    4624: romdata_int <= 'h1706;
    4625: romdata_int <= 'h240b;
    4626: romdata_int <= 'h67b;
    4627: romdata_int <= 'h203e;
    4628: romdata_int <= 'h1edb;
    4629: romdata_int <= 'h2958;
    4630: romdata_int <= 'h8ee;
    4631: romdata_int <= 'h28c3;
    4632: romdata_int <= 'h1c45;
    4633: romdata_int <= 'h487;
    4634: romdata_int <= 'h285c;
    4635: romdata_int <= 'h181e; // Line Descriptor
    4636: romdata_int <= 'hc00;
    4637: romdata_int <= 'h2282;
    4638: romdata_int <= 'h2a67;
    4639: romdata_int <= 'h3473;
    4640: romdata_int <= 'h1c2b;
    4641: romdata_int <= 'h1758;
    4642: romdata_int <= 'h3ac5;
    4643: romdata_int <= 'h12ad;
    4644: romdata_int <= 'h2a35;
    4645: romdata_int <= 'h1642;
    4646: romdata_int <= 'h1217;
    4647: romdata_int <= 'hd15;
    4648: romdata_int <= 'h14c;
    4649: romdata_int <= 'h181e; // Line Descriptor
    4650: romdata_int <= 'he00;
    4651: romdata_int <= 'h1ae5;
    4652: romdata_int <= 'h366b;
    4653: romdata_int <= 'he39;
    4654: romdata_int <= 'h1966;
    4655: romdata_int <= 'h307;
    4656: romdata_int <= 'h1d45;
    4657: romdata_int <= 'ha9e;
    4658: romdata_int <= 'h2481;
    4659: romdata_int <= 'h274d;
    4660: romdata_int <= 'hc8b;
    4661: romdata_int <= 'h3099;
    4662: romdata_int <= 'he34;
    4663: romdata_int <= 'h181e; // Line Descriptor
    4664: romdata_int <= 'h1000;
    4665: romdata_int <= 'h3760;
    4666: romdata_int <= 'ha49;
    4667: romdata_int <= 'h1238;
    4668: romdata_int <= 'h3862;
    4669: romdata_int <= 'h28b4;
    4670: romdata_int <= 'h56;
    4671: romdata_int <= 'h660;
    4672: romdata_int <= 'h20d8;
    4673: romdata_int <= 'h2a03;
    4674: romdata_int <= 'h2ec8;
    4675: romdata_int <= 'h822;
    4676: romdata_int <= 'h1294;
    4677: romdata_int <= 'h181e; // Line Descriptor
    4678: romdata_int <= 'h1200;
    4679: romdata_int <= 'hc7e;
    4680: romdata_int <= 'h1b1e;
    4681: romdata_int <= 'h845;
    4682: romdata_int <= 'h2a6e;
    4683: romdata_int <= 'h22a8;
    4684: romdata_int <= 'h1430;
    4685: romdata_int <= 'h80;
    4686: romdata_int <= 'h1cb5;
    4687: romdata_int <= 'h4db;
    4688: romdata_int <= 'h867;
    4689: romdata_int <= 'h2d49;
    4690: romdata_int <= 'h1832;
    4691: romdata_int <= 'h181e; // Line Descriptor
    4692: romdata_int <= 'h1400;
    4693: romdata_int <= 'h391c;
    4694: romdata_int <= 'h243d;
    4695: romdata_int <= 'h2d59;
    4696: romdata_int <= 'h3298;
    4697: romdata_int <= 'h2ef3;
    4698: romdata_int <= 'h34d9;
    4699: romdata_int <= 'h26d4;
    4700: romdata_int <= 'h343a;
    4701: romdata_int <= 'h193b;
    4702: romdata_int <= 'h3451;
    4703: romdata_int <= 'h34ba;
    4704: romdata_int <= 'h1f4c;
    4705: romdata_int <= 'h181e; // Line Descriptor
    4706: romdata_int <= 'h1600;
    4707: romdata_int <= 'h1d11;
    4708: romdata_int <= 'h761;
    4709: romdata_int <= 'h1f08;
    4710: romdata_int <= 'hc79;
    4711: romdata_int <= 'h1881;
    4712: romdata_int <= 'h80d;
    4713: romdata_int <= 'h38c6;
    4714: romdata_int <= 'h171d;
    4715: romdata_int <= 'h324f;
    4716: romdata_int <= 'h3af2;
    4717: romdata_int <= 'h3734;
    4718: romdata_int <= 'h254c;
    4719: romdata_int <= 'h181e; // Line Descriptor
    4720: romdata_int <= 'h1800;
    4721: romdata_int <= 'h3303;
    4722: romdata_int <= 'h1c02;
    4723: romdata_int <= 'h1a36;
    4724: romdata_int <= 'h53e;
    4725: romdata_int <= 'h36e4;
    4726: romdata_int <= 'h4f5;
    4727: romdata_int <= 'h36d5;
    4728: romdata_int <= 'h10fc;
    4729: romdata_int <= 'h762;
    4730: romdata_int <= 'ha18;
    4731: romdata_int <= 'h1654;
    4732: romdata_int <= 'h332f;
    4733: romdata_int <= 'h181e; // Line Descriptor
    4734: romdata_int <= 'h1a00;
    4735: romdata_int <= 'h16ee;
    4736: romdata_int <= 'h2c52;
    4737: romdata_int <= 'h8e;
    4738: romdata_int <= 'h2ea6;
    4739: romdata_int <= 'h3350;
    4740: romdata_int <= 'h12f7;
    4741: romdata_int <= 'h2f32;
    4742: romdata_int <= 'h2df;
    4743: romdata_int <= 'h1125;
    4744: romdata_int <= 'h2c45;
    4745: romdata_int <= 'h1b13;
    4746: romdata_int <= 'ha7d;
    4747: romdata_int <= 'h181e; // Line Descriptor
    4748: romdata_int <= 'h1c00;
    4749: romdata_int <= 'h78;
    4750: romdata_int <= 'h13;
    4751: romdata_int <= 'h3696;
    4752: romdata_int <= 'h2806;
    4753: romdata_int <= 'h3943;
    4754: romdata_int <= 'h2ae1;
    4755: romdata_int <= 'h1e42;
    4756: romdata_int <= 'h2d28;
    4757: romdata_int <= 'h20b5;
    4758: romdata_int <= 'h2419;
    4759: romdata_int <= 'h2e24;
    4760: romdata_int <= 'h14d9;
    4761: romdata_int <= 'h41e; // Line Descriptor
    4762: romdata_int <= 'h1e00;
    4763: romdata_int <= 'h8d2;
    4764: romdata_int <= 'h2fe;
    4765: romdata_int <= 'h41e; // Line Descriptor
    4766: romdata_int <= 'h2000;
    4767: romdata_int <= 'h24d8;
    4768: romdata_int <= 'h3b32;
    4769: romdata_int <= 'h41e; // Line Descriptor
    4770: romdata_int <= 'h2200;
    4771: romdata_int <= 'h6f3;
    4772: romdata_int <= 'hce2;
    4773: romdata_int <= 'h41e; // Line Descriptor
    4774: romdata_int <= 'h2400;
    4775: romdata_int <= 'h14c6;
    4776: romdata_int <= 'h3838;
    4777: romdata_int <= 'h41e; // Line Descriptor
    4778: romdata_int <= 'h2600;
    4779: romdata_int <= 'h31c;
    4780: romdata_int <= 'h2e3b;
    4781: romdata_int <= 'h41e; // Line Descriptor
    4782: romdata_int <= 'h2800;
    4783: romdata_int <= 'h30cd;
    4784: romdata_int <= 'h3105;
    4785: romdata_int <= 'h41e; // Line Descriptor
    4786: romdata_int <= 'h2a00;
    4787: romdata_int <= 'h2f45;
    4788: romdata_int <= 'h2827;
    4789: romdata_int <= 'h41e; // Line Descriptor
    4790: romdata_int <= 'h2c00;
    4791: romdata_int <= 'hf3d;
    4792: romdata_int <= 'h1156;
    4793: romdata_int <= 'h41e; // Line Descriptor
    4794: romdata_int <= 'h2e00;
    4795: romdata_int <= 'h2a48;
    4796: romdata_int <= 'h2737;
    4797: romdata_int <= 'h41e; // Line Descriptor
    4798: romdata_int <= 'h3000;
    4799: romdata_int <= 'h3a40;
    4800: romdata_int <= 'h14b9;
    4801: romdata_int <= 'h41e; // Line Descriptor
    4802: romdata_int <= 'h3200;
    4803: romdata_int <= 'h3433;
    4804: romdata_int <= 'h1e12;
    4805: romdata_int <= 'h41e; // Line Descriptor
    4806: romdata_int <= 'h3400;
    4807: romdata_int <= 'h291e;
    4808: romdata_int <= 'h227f;
    4809: romdata_int <= 'h41e; // Line Descriptor
    4810: romdata_int <= 'h3600;
    4811: romdata_int <= 'h4a9;
    4812: romdata_int <= 'he23;
    4813: romdata_int <= 'h41e; // Line Descriptor
    4814: romdata_int <= 'h3800;
    4815: romdata_int <= 'h1108;
    4816: romdata_int <= 'h476;
    4817: romdata_int <= 'h41e; // Line Descriptor
    4818: romdata_int <= 'h3a00;
    4819: romdata_int <= 'h206b;
    4820: romdata_int <= 'h187d;
    4821: romdata_int <= 'h41e; // Line Descriptor
    4822: romdata_int <= 'h0;
    4823: romdata_int <= 'h32ea;
    4824: romdata_int <= 'h2850;
    4825: romdata_int <= 'h41e; // Line Descriptor
    4826: romdata_int <= 'h200;
    4827: romdata_int <= 'h1f41;
    4828: romdata_int <= 'h258;
    4829: romdata_int <= 'h41e; // Line Descriptor
    4830: romdata_int <= 'h400;
    4831: romdata_int <= 'h1c5c;
    4832: romdata_int <= 'h2c51;
    4833: romdata_int <= 'h41e; // Line Descriptor
    4834: romdata_int <= 'h600;
    4835: romdata_int <= 'h2ab1;
    4836: romdata_int <= 'h2a43;
    4837: romdata_int <= 'h41e; // Line Descriptor
    4838: romdata_int <= 'h800;
    4839: romdata_int <= 'h1539;
    4840: romdata_int <= 'h6fa;
    4841: romdata_int <= 'h41e; // Line Descriptor
    4842: romdata_int <= 'ha00;
    4843: romdata_int <= 'h283d;
    4844: romdata_int <= 'h384d;
    4845: romdata_int <= 'h41e; // Line Descriptor
    4846: romdata_int <= 'hc00;
    4847: romdata_int <= 'h215c;
    4848: romdata_int <= 'h3145;
    4849: romdata_int <= 'h41e; // Line Descriptor
    4850: romdata_int <= 'he00;
    4851: romdata_int <= 'h1838;
    4852: romdata_int <= 'hd35;
    4853: romdata_int <= 'h41e; // Line Descriptor
    4854: romdata_int <= 'h1000;
    4855: romdata_int <= 'h234e;
    4856: romdata_int <= 'h2486;
    4857: romdata_int <= 'h41e; // Line Descriptor
    4858: romdata_int <= 'h1200;
    4859: romdata_int <= 'h884;
    4860: romdata_int <= 'h100b;
    4861: romdata_int <= 'h41e; // Line Descriptor
    4862: romdata_int <= 'h1400;
    4863: romdata_int <= 'h58;
    4864: romdata_int <= 'h22a9;
    4865: romdata_int <= 'h41e; // Line Descriptor
    4866: romdata_int <= 'h1600;
    4867: romdata_int <= 'h241c;
    4868: romdata_int <= 'h2e73;
    4869: romdata_int <= 'h41e; // Line Descriptor
    4870: romdata_int <= 'h1800;
    4871: romdata_int <= 'h4ba;
    4872: romdata_int <= 'h1abd;
    4873: romdata_int <= 'h41e; // Line Descriptor
    4874: romdata_int <= 'h1a00;
    4875: romdata_int <= 'h1b3d;
    4876: romdata_int <= 'h201e;
    4877: romdata_int <= 'h41e; // Line Descriptor
    4878: romdata_int <= 'h1c00;
    4879: romdata_int <= 'h3688;
    4880: romdata_int <= 'h3a33;
    4881: romdata_int <= 'h41e; // Line Descriptor
    4882: romdata_int <= 'h1e00;
    4883: romdata_int <= 'hc96;
    4884: romdata_int <= 'h1674;
    4885: romdata_int <= 'h41e; // Line Descriptor
    4886: romdata_int <= 'h2000;
    4887: romdata_int <= 'h311;
    4888: romdata_int <= 'h188b;
    4889: romdata_int <= 'h41e; // Line Descriptor
    4890: romdata_int <= 'h2200;
    4891: romdata_int <= 'h2d53;
    4892: romdata_int <= 'hecd;
    4893: romdata_int <= 'h41e; // Line Descriptor
    4894: romdata_int <= 'h2400;
    4895: romdata_int <= 'h38bc;
    4896: romdata_int <= 'ha6e;
    4897: romdata_int <= 'h41e; // Line Descriptor
    4898: romdata_int <= 'h2600;
    4899: romdata_int <= 'h3a72;
    4900: romdata_int <= 'h1433;
    4901: romdata_int <= 'h41e; // Line Descriptor
    4902: romdata_int <= 'h2800;
    4903: romdata_int <= 'h349e;
    4904: romdata_int <= 'h3659;
    4905: romdata_int <= 'h41e; // Line Descriptor
    4906: romdata_int <= 'h2a00;
    4907: romdata_int <= 'h2687;
    4908: romdata_int <= 'h1ede;
    4909: romdata_int <= 'h41e; // Line Descriptor
    4910: romdata_int <= 'h2c00;
    4911: romdata_int <= 'he25;
    4912: romdata_int <= 'h3421;
    4913: romdata_int <= 'h41e; // Line Descriptor
    4914: romdata_int <= 'h2e00;
    4915: romdata_int <= 'h12bb;
    4916: romdata_int <= 'h3266;
    4917: romdata_int <= 'h41e; // Line Descriptor
    4918: romdata_int <= 'h3000;
    4919: romdata_int <= 'h2f1a;
    4920: romdata_int <= 'h118;
    4921: romdata_int <= 'h41e; // Line Descriptor
    4922: romdata_int <= 'h3200;
    4923: romdata_int <= 'hb13;
    4924: romdata_int <= 'h80d;
    4925: romdata_int <= 'h41e; // Line Descriptor
    4926: romdata_int <= 'h3400;
    4927: romdata_int <= 'h10d3;
    4928: romdata_int <= 'h4a8;
    4929: romdata_int <= 'h41e; // Line Descriptor
    4930: romdata_int <= 'h3600;
    4931: romdata_int <= 'h30cd;
    4932: romdata_int <= 'h26aa;
    4933: romdata_int <= 'h41e; // Line Descriptor
    4934: romdata_int <= 'h3800;
    4935: romdata_int <= 'h6f0;
    4936: romdata_int <= 'h1242;
    4937: romdata_int <= 'h41e; // Line Descriptor
    4938: romdata_int <= 'h3a00;
    4939: romdata_int <= 'h163b;
    4940: romdata_int <= 'h1cac;
    4941: romdata_int <= 'h41e; // Line Descriptor
    4942: romdata_int <= 'h0;
    4943: romdata_int <= 'h3030;
    4944: romdata_int <= 'h2676;
    4945: romdata_int <= 'h41e; // Line Descriptor
    4946: romdata_int <= 'h200;
    4947: romdata_int <= 'h2070;
    4948: romdata_int <= 'h1c8c;
    4949: romdata_int <= 'h41e; // Line Descriptor
    4950: romdata_int <= 'h400;
    4951: romdata_int <= 'h10f1;
    4952: romdata_int <= 'he02;
    4953: romdata_int <= 'h41e; // Line Descriptor
    4954: romdata_int <= 'h600;
    4955: romdata_int <= 'hb61;
    4956: romdata_int <= 'h1726;
    4957: romdata_int <= 'h41e; // Line Descriptor
    4958: romdata_int <= 'h800;
    4959: romdata_int <= 'h2a28;
    4960: romdata_int <= 'h6d9;
    4961: romdata_int <= 'h41e; // Line Descriptor
    4962: romdata_int <= 'ha00;
    4963: romdata_int <= 'h28b0;
    4964: romdata_int <= 'h49b;
    4965: romdata_int <= 'h41e; // Line Descriptor
    4966: romdata_int <= 'hc00;
    4967: romdata_int <= 'h262f;
    4968: romdata_int <= 'h3b44;
    4969: romdata_int <= 'h41e; // Line Descriptor
    4970: romdata_int <= 'he00;
    4971: romdata_int <= 'h2506;
    4972: romdata_int <= 'h2ab;
    4973: romdata_int <= 'h41e; // Line Descriptor
    4974: romdata_int <= 'h1000;
    4975: romdata_int <= 'h3293;
    4976: romdata_int <= 'h3156;
    4977: romdata_int <= 'h41e; // Line Descriptor
    4978: romdata_int <= 'h1200;
    4979: romdata_int <= 'h2d3;
    4980: romdata_int <= 'h22b7;
    4981: romdata_int <= 'h41e; // Line Descriptor
    4982: romdata_int <= 'h1400;
    4983: romdata_int <= 'h4de;
    4984: romdata_int <= 'h2aa4;
    4985: romdata_int <= 'h41e; // Line Descriptor
    4986: romdata_int <= 'h1600;
    4987: romdata_int <= 'h1d40;
    4988: romdata_int <= 'h1155;
    4989: romdata_int <= 'h41e; // Line Descriptor
    4990: romdata_int <= 'h1800;
    4991: romdata_int <= 'h118;
    4992: romdata_int <= 'h1f0b;
    4993: romdata_int <= 'h41e; // Line Descriptor
    4994: romdata_int <= 'h1a00;
    4995: romdata_int <= 'hd31;
    4996: romdata_int <= 'h28bb;
    4997: romdata_int <= 'h41e; // Line Descriptor
    4998: romdata_int <= 'h1c00;
    4999: romdata_int <= 'h22eb;
    5000: romdata_int <= 'h3927;
    5001: romdata_int <= 'h41e; // Line Descriptor
    5002: romdata_int <= 'h1e00;
    5003: romdata_int <= 'h372c;
    5004: romdata_int <= 'h3271;
    5005: romdata_int <= 'h41e; // Line Descriptor
    5006: romdata_int <= 'h2000;
    5007: romdata_int <= 'h1438;
    5008: romdata_int <= 'h3480;
    5009: romdata_int <= 'h41e; // Line Descriptor
    5010: romdata_int <= 'h2200;
    5011: romdata_int <= 'h85f;
    5012: romdata_int <= 'h131a;
    5013: romdata_int <= 'h41e; // Line Descriptor
    5014: romdata_int <= 'h2400;
    5015: romdata_int <= 'h34ce;
    5016: romdata_int <= 'h15;
    5017: romdata_int <= 'h41e; // Line Descriptor
    5018: romdata_int <= 'h2600;
    5019: romdata_int <= 'h60c;
    5020: romdata_int <= 'h2eb5;
    5021: romdata_int <= 'h41e; // Line Descriptor
    5022: romdata_int <= 'h2800;
    5023: romdata_int <= 'h1e89;
    5024: romdata_int <= 'h24e9;
    5025: romdata_int <= 'h41e; // Line Descriptor
    5026: romdata_int <= 'h2a00;
    5027: romdata_int <= 'h2c35;
    5028: romdata_int <= 'h18df;
    5029: romdata_int <= 'h41e; // Line Descriptor
    5030: romdata_int <= 'h2c00;
    5031: romdata_int <= 'h132e;
    5032: romdata_int <= 'h2133;
    5033: romdata_int <= 'h41e; // Line Descriptor
    5034: romdata_int <= 'h2e00;
    5035: romdata_int <= 'hec0;
    5036: romdata_int <= 'h1487;
    5037: romdata_int <= 'h41e; // Line Descriptor
    5038: romdata_int <= 'h3000;
    5039: romdata_int <= 'h2e7c;
    5040: romdata_int <= 'h3733;
    5041: romdata_int <= 'h41e; // Line Descriptor
    5042: romdata_int <= 'h3200;
    5043: romdata_int <= 'h38e9;
    5044: romdata_int <= 'h2cb9;
    5045: romdata_int <= 'h41e; // Line Descriptor
    5046: romdata_int <= 'h3400;
    5047: romdata_int <= 'h1928;
    5048: romdata_int <= 'hc97;
    5049: romdata_int <= 'h41e; // Line Descriptor
    5050: romdata_int <= 'h3600;
    5051: romdata_int <= 'h1a1c;
    5052: romdata_int <= 'h8ca;
    5053: romdata_int <= 'h41e; // Line Descriptor
    5054: romdata_int <= 'h3800;
    5055: romdata_int <= 'h3b0c;
    5056: romdata_int <= 'h1ac4;
    5057: romdata_int <= 'h41e; // Line Descriptor
    5058: romdata_int <= 'h3a00;
    5059: romdata_int <= 'h1644;
    5060: romdata_int <= 'ha60;
    5061: romdata_int <= 'h41e; // Line Descriptor
    5062: romdata_int <= 'h0;
    5063: romdata_int <= 'h1764;
    5064: romdata_int <= 'h669;
    5065: romdata_int <= 'h41e; // Line Descriptor
    5066: romdata_int <= 'h200;
    5067: romdata_int <= 'h478;
    5068: romdata_int <= 'ha87;
    5069: romdata_int <= 'h41e; // Line Descriptor
    5070: romdata_int <= 'h400;
    5071: romdata_int <= 'h380a;
    5072: romdata_int <= 'he39;
    5073: romdata_int <= 'h41e; // Line Descriptor
    5074: romdata_int <= 'h600;
    5075: romdata_int <= 'h3a49;
    5076: romdata_int <= 'h3b35;
    5077: romdata_int <= 'h41e; // Line Descriptor
    5078: romdata_int <= 'h800;
    5079: romdata_int <= 'h2640;
    5080: romdata_int <= 'h1107;
    5081: romdata_int <= 'h41e; // Line Descriptor
    5082: romdata_int <= 'ha00;
    5083: romdata_int <= 'h2214;
    5084: romdata_int <= 'h3406;
    5085: romdata_int <= 'h41e; // Line Descriptor
    5086: romdata_int <= 'hc00;
    5087: romdata_int <= 'h311c;
    5088: romdata_int <= 'h302d;
    5089: romdata_int <= 'h41e; // Line Descriptor
    5090: romdata_int <= 'he00;
    5091: romdata_int <= 'h3563;
    5092: romdata_int <= 'h6c;
    5093: romdata_int <= 'h41e; // Line Descriptor
    5094: romdata_int <= 'h1000;
    5095: romdata_int <= 'h18de;
    5096: romdata_int <= 'h133c;
    5097: romdata_int <= 'h41e; // Line Descriptor
    5098: romdata_int <= 'h1200;
    5099: romdata_int <= 'h2869;
    5100: romdata_int <= 'h22f8;
    5101: romdata_int <= 'h41e; // Line Descriptor
    5102: romdata_int <= 'h1400;
    5103: romdata_int <= 'h1106;
    5104: romdata_int <= 'h2bf;
    5105: romdata_int <= 'h41e; // Line Descriptor
    5106: romdata_int <= 'h1600;
    5107: romdata_int <= 'h2cc;
    5108: romdata_int <= 'h2d65;
    5109: romdata_int <= 'h41e; // Line Descriptor
    5110: romdata_int <= 'h1800;
    5111: romdata_int <= 'h1aa1;
    5112: romdata_int <= 'h1930;
    5113: romdata_int <= 'h41e; // Line Descriptor
    5114: romdata_int <= 'h1a00;
    5115: romdata_int <= 'h1413;
    5116: romdata_int <= 'h2b3f;
    5117: romdata_int <= 'h41e; // Line Descriptor
    5118: romdata_int <= 'h1c00;
    5119: romdata_int <= 'h36d0;
    5120: romdata_int <= 'h2935;
    5121: romdata_int <= 'h41e; // Line Descriptor
    5122: romdata_int <= 'h1e00;
    5123: romdata_int <= 'h1264;
    5124: romdata_int <= 'h244b;
    5125: romdata_int <= 'h41e; // Line Descriptor
    5126: romdata_int <= 'h2000;
    5127: romdata_int <= 'h1e06;
    5128: romdata_int <= 'h2650;
    5129: romdata_int <= 'h41e; // Line Descriptor
    5130: romdata_int <= 'h2200;
    5131: romdata_int <= 'hd0b;
    5132: romdata_int <= 'h3633;
    5133: romdata_int <= 'h41e; // Line Descriptor
    5134: romdata_int <= 'h2400;
    5135: romdata_int <= 'h2032;
    5136: romdata_int <= 'h1f32;
    5137: romdata_int <= 'h41e; // Line Descriptor
    5138: romdata_int <= 'h2600;
    5139: romdata_int <= 'h2d0c;
    5140: romdata_int <= 'h92e;
    5141: romdata_int <= 'h41e; // Line Descriptor
    5142: romdata_int <= 'h2800;
    5143: romdata_int <= 'h3245;
    5144: romdata_int <= 'h392a;
    5145: romdata_int <= 'h41e; // Line Descriptor
    5146: romdata_int <= 'h2a00;
    5147: romdata_int <= 'h619;
    5148: romdata_int <= 'hcf4;
    5149: romdata_int <= 'h41e; // Line Descriptor
    5150: romdata_int <= 'h2c00;
    5151: romdata_int <= 'h2ad1;
    5152: romdata_int <= 'h2e7f;
    5153: romdata_int <= 'h41e; // Line Descriptor
    5154: romdata_int <= 'h2e00;
    5155: romdata_int <= 'h857;
    5156: romdata_int <= 'h1d05;
    5157: romdata_int <= 'h41e; // Line Descriptor
    5158: romdata_int <= 'h3000;
    5159: romdata_int <= 'h2e4c;
    5160: romdata_int <= 'h2015;
    5161: romdata_int <= 'h41e; // Line Descriptor
    5162: romdata_int <= 'h3200;
    5163: romdata_int <= 'ha45;
    5164: romdata_int <= 'h1614;
    5165: romdata_int <= 'h41e; // Line Descriptor
    5166: romdata_int <= 'h3400;
    5167: romdata_int <= 'he9c;
    5168: romdata_int <= 'h40c;
    5169: romdata_int <= 'h41e; // Line Descriptor
    5170: romdata_int <= 'h3600;
    5171: romdata_int <= 'h1d21;
    5172: romdata_int <= 'h154b;
    5173: romdata_int <= 'h41e; // Line Descriptor
    5174: romdata_int <= 'h3800;
    5175: romdata_int <= 'ha1;
    5176: romdata_int <= 'h3244;
    5177: romdata_int <= 'h41e; // Line Descriptor
    5178: romdata_int <= 'h3a00;
    5179: romdata_int <= 'h24ea;
    5180: romdata_int <= 'h1a2d;
    5181: romdata_int <= 'h41e; // Line Descriptor
    5182: romdata_int <= 'h0;
    5183: romdata_int <= 'h3a3a;
    5184: romdata_int <= 'hf05;
    5185: romdata_int <= 'h41e; // Line Descriptor
    5186: romdata_int <= 'h200;
    5187: romdata_int <= 'h2a7e;
    5188: romdata_int <= 'h1238;
    5189: romdata_int <= 'h41e; // Line Descriptor
    5190: romdata_int <= 'h400;
    5191: romdata_int <= 'h294f;
    5192: romdata_int <= 'h264e;
    5193: romdata_int <= 'h41e; // Line Descriptor
    5194: romdata_int <= 'h600;
    5195: romdata_int <= 'he7a;
    5196: romdata_int <= 'h254a;
    5197: romdata_int <= 'h41e; // Line Descriptor
    5198: romdata_int <= 'h800;
    5199: romdata_int <= 'h303f;
    5200: romdata_int <= 'h28e6;
    5201: romdata_int <= 'h41e; // Line Descriptor
    5202: romdata_int <= 'ha00;
    5203: romdata_int <= 'h1c8d;
    5204: romdata_int <= 'h3abc;
    5205: romdata_int <= 'h41e; // Line Descriptor
    5206: romdata_int <= 'hc00;
    5207: romdata_int <= 'h1f55;
    5208: romdata_int <= 'h2b04;
    5209: romdata_int <= 'h41e; // Line Descriptor
    5210: romdata_int <= 'he00;
    5211: romdata_int <= 'h38fe;
    5212: romdata_int <= 'h1c83;
    5213: romdata_int <= 'h41e; // Line Descriptor
    5214: romdata_int <= 'h1000;
    5215: romdata_int <= 'h146e;
    5216: romdata_int <= 'h38b6;
    5217: romdata_int <= 'h41e; // Line Descriptor
    5218: romdata_int <= 'h1200;
    5219: romdata_int <= 'h20d3;
    5220: romdata_int <= 'hd42;
    5221: romdata_int <= 'h41e; // Line Descriptor
    5222: romdata_int <= 'h1400;
    5223: romdata_int <= 'h10ec;
    5224: romdata_int <= 'h4cc;
    5225: romdata_int <= 'h41e; // Line Descriptor
    5226: romdata_int <= 'h1600;
    5227: romdata_int <= 'h22b;
    5228: romdata_int <= 'h3704;
    5229: romdata_int <= 'h41e; // Line Descriptor
    5230: romdata_int <= 'h1800;
    5231: romdata_int <= 'h561;
    5232: romdata_int <= 'hb2a;
    5233: romdata_int <= 'h41e; // Line Descriptor
    5234: romdata_int <= 'h1a00;
    5235: romdata_int <= 'h1278;
    5236: romdata_int <= 'h14ed;
    5237: romdata_int <= 'h41e; // Line Descriptor
    5238: romdata_int <= 'h1c00;
    5239: romdata_int <= 'h2531;
    5240: romdata_int <= 'h2d2f;
    5241: romdata_int <= 'h41e; // Line Descriptor
    5242: romdata_int <= 'h1e00;
    5243: romdata_int <= 'h2ece;
    5244: romdata_int <= 'h190c;
    5245: romdata_int <= 'h41e; // Line Descriptor
    5246: romdata_int <= 'h2000;
    5247: romdata_int <= 'h6f;
    5248: romdata_int <= 'h1e60;
    5249: romdata_int <= 'h41e; // Line Descriptor
    5250: romdata_int <= 'h2200;
    5251: romdata_int <= 'h88e;
    5252: romdata_int <= 'h760;
    5253: romdata_int <= 'h41e; // Line Descriptor
    5254: romdata_int <= 'h2400;
    5255: romdata_int <= 'h355f;
    5256: romdata_int <= 'h20d8;
    5257: romdata_int <= 'h41e; // Line Descriptor
    5258: romdata_int <= 'h2600;
    5259: romdata_int <= 'h2325;
    5260: romdata_int <= 'h32fe;
    5261: romdata_int <= 'h41e; // Line Descriptor
    5262: romdata_int <= 'h2800;
    5263: romdata_int <= 'h2642;
    5264: romdata_int <= 'h97;
    5265: romdata_int <= 'h41e; // Line Descriptor
    5266: romdata_int <= 'h2a00;
    5267: romdata_int <= 'h2d32;
    5268: romdata_int <= 'h10e3;
    5269: romdata_int <= 'h41e; // Line Descriptor
    5270: romdata_int <= 'h2c00;
    5271: romdata_int <= 'h1a71;
    5272: romdata_int <= 'h3039;
    5273: romdata_int <= 'h41e; // Line Descriptor
    5274: romdata_int <= 'h2e00;
    5275: romdata_int <= 'hc46;
    5276: romdata_int <= 'h2f2c;
    5277: romdata_int <= 'h41e; // Line Descriptor
    5278: romdata_int <= 'h3000;
    5279: romdata_int <= 'h16e5;
    5280: romdata_int <= 'h1a81;
    5281: romdata_int <= 'h41e; // Line Descriptor
    5282: romdata_int <= 'h3200;
    5283: romdata_int <= 'h3281;
    5284: romdata_int <= 'h1648;
    5285: romdata_int <= 'h41e; // Line Descriptor
    5286: romdata_int <= 'h3400;
    5287: romdata_int <= 'h1887;
    5288: romdata_int <= 'h8d6;
    5289: romdata_int <= 'h41e; // Line Descriptor
    5290: romdata_int <= 'h3600;
    5291: romdata_int <= 'ha7d;
    5292: romdata_int <= 'h353d;
    5293: romdata_int <= 'h41e; // Line Descriptor
    5294: romdata_int <= 'h3800;
    5295: romdata_int <= 'h69c;
    5296: romdata_int <= 'h247;
    5297: romdata_int <= 'h51e; // Line Descriptor
    5298: romdata_int <= 'h3a00;
    5299: romdata_int <= 'h36f4;
    5300: romdata_int <= 'h230b;
    5301: romdata_int <= 'h614; // Line Descriptor
    5302: romdata_int <= 'h0;
    5303: romdata_int <= 'h1f37;
    5304: romdata_int <= 'h108e;
    5305: romdata_int <= 'h4a1;
    5306: romdata_int <= 'h614; // Line Descriptor
    5307: romdata_int <= 'h200;
    5308: romdata_int <= 'h122;
    5309: romdata_int <= 'h18ae;
    5310: romdata_int <= 'h110b;
    5311: romdata_int <= 'h614; // Line Descriptor
    5312: romdata_int <= 'h400;
    5313: romdata_int <= 'h2289;
    5314: romdata_int <= 'he2e;
    5315: romdata_int <= 'h1404;
    5316: romdata_int <= 'h614; // Line Descriptor
    5317: romdata_int <= 'h600;
    5318: romdata_int <= 'h35c;
    5319: romdata_int <= 'h20e1;
    5320: romdata_int <= 'h26ec;
    5321: romdata_int <= 'h614; // Line Descriptor
    5322: romdata_int <= 'h800;
    5323: romdata_int <= 'h183a;
    5324: romdata_int <= 'h22a1;
    5325: romdata_int <= 'h939;
    5326: romdata_int <= 'h614; // Line Descriptor
    5327: romdata_int <= 'ha00;
    5328: romdata_int <= 'he60;
    5329: romdata_int <= 'ha79;
    5330: romdata_int <= 'h6b8;
    5331: romdata_int <= 'h614; // Line Descriptor
    5332: romdata_int <= 'hc00;
    5333: romdata_int <= 'h1cb9;
    5334: romdata_int <= 'h133b;
    5335: romdata_int <= 'h1e7c;
    5336: romdata_int <= 'h614; // Line Descriptor
    5337: romdata_int <= 'he00;
    5338: romdata_int <= 'h1499;
    5339: romdata_int <= 'h53d;
    5340: romdata_int <= 'h1d65;
    5341: romdata_int <= 'h614; // Line Descriptor
    5342: romdata_int <= 'h1000;
    5343: romdata_int <= 'h1079;
    5344: romdata_int <= 'h1a1e;
    5345: romdata_int <= 'h2bc;
    5346: romdata_int <= 'h614; // Line Descriptor
    5347: romdata_int <= 'h1200;
    5348: romdata_int <= 'hc91;
    5349: romdata_int <= 'h80d;
    5350: romdata_int <= 'hf28;
    5351: romdata_int <= 'h614; // Line Descriptor
    5352: romdata_int <= 'h1400;
    5353: romdata_int <= 'h2055;
    5354: romdata_int <= 'h1461;
    5355: romdata_int <= 'h1ad5;
    5356: romdata_int <= 'h614; // Line Descriptor
    5357: romdata_int <= 'h1600;
    5358: romdata_int <= 'h1ae6;
    5359: romdata_int <= 'h2734;
    5360: romdata_int <= 'h16ae;
    5361: romdata_int <= 'h614; // Line Descriptor
    5362: romdata_int <= 'h1800;
    5363: romdata_int <= 'haf3;
    5364: romdata_int <= 'hca4;
    5365: romdata_int <= 'hb2c;
    5366: romdata_int <= 'h614; // Line Descriptor
    5367: romdata_int <= 'h1a00;
    5368: romdata_int <= 'h643;
    5369: romdata_int <= 'h728;
    5370: romdata_int <= 'h12b0;
    5371: romdata_int <= 'h614; // Line Descriptor
    5372: romdata_int <= 'h1c00;
    5373: romdata_int <= 'h12e5;
    5374: romdata_int <= 'h1ec9;
    5375: romdata_int <= 'h186a;
    5376: romdata_int <= 'h614; // Line Descriptor
    5377: romdata_int <= 'h1e00;
    5378: romdata_int <= 'h264e;
    5379: romdata_int <= 'hc4;
    5380: romdata_int <= 'h2350;
    5381: romdata_int <= 'h614; // Line Descriptor
    5382: romdata_int <= 'h2000;
    5383: romdata_int <= 'h852;
    5384: romdata_int <= 'h163b;
    5385: romdata_int <= 'h252b;
    5386: romdata_int <= 'h614; // Line Descriptor
    5387: romdata_int <= 'h2200;
    5388: romdata_int <= 'h44a;
    5389: romdata_int <= 'h277;
    5390: romdata_int <= 'he7;
    5391: romdata_int <= 'h614; // Line Descriptor
    5392: romdata_int <= 'h2400;
    5393: romdata_int <= 'h1753;
    5394: romdata_int <= 'h1d2c;
    5395: romdata_int <= 'h2149;
    5396: romdata_int <= 'h614; // Line Descriptor
    5397: romdata_int <= 'h2600;
    5398: romdata_int <= 'h2488;
    5399: romdata_int <= 'h2527;
    5400: romdata_int <= 'hcbd;
    5401: romdata_int <= 'h414; // Line Descriptor
    5402: romdata_int <= 'h0;
    5403: romdata_int <= 'h2101;
    5404: romdata_int <= 'hd34;
    5405: romdata_int <= 'h414; // Line Descriptor
    5406: romdata_int <= 'h200;
    5407: romdata_int <= 'h84b;
    5408: romdata_int <= 'h20d9;
    5409: romdata_int <= 'h414; // Line Descriptor
    5410: romdata_int <= 'h400;
    5411: romdata_int <= 'h1406;
    5412: romdata_int <= 'h85f;
    5413: romdata_int <= 'h414; // Line Descriptor
    5414: romdata_int <= 'h600;
    5415: romdata_int <= 'hf2d;
    5416: romdata_int <= 'he9f;
    5417: romdata_int <= 'h414; // Line Descriptor
    5418: romdata_int <= 'h800;
    5419: romdata_int <= 'h254f;
    5420: romdata_int <= 'h2625;
    5421: romdata_int <= 'h414; // Line Descriptor
    5422: romdata_int <= 'ha00;
    5423: romdata_int <= 'h138;
    5424: romdata_int <= 'h148f;
    5425: romdata_int <= 'h414; // Line Descriptor
    5426: romdata_int <= 'hc00;
    5427: romdata_int <= 'h675;
    5428: romdata_int <= 'h1641;
    5429: romdata_int <= 'h414; // Line Descriptor
    5430: romdata_int <= 'he00;
    5431: romdata_int <= 'h2633;
    5432: romdata_int <= 'hb11;
    5433: romdata_int <= 'h414; // Line Descriptor
    5434: romdata_int <= 'h1000;
    5435: romdata_int <= 'h234a;
    5436: romdata_int <= 'h1a7d;
    5437: romdata_int <= 'h414; // Line Descriptor
    5438: romdata_int <= 'h1200;
    5439: romdata_int <= 'h104f;
    5440: romdata_int <= 'h505;
    5441: romdata_int <= 'h414; // Line Descriptor
    5442: romdata_int <= 'h1400;
    5443: romdata_int <= 'h348;
    5444: romdata_int <= 'h1e1a;
    5445: romdata_int <= 'h414; // Line Descriptor
    5446: romdata_int <= 'h1600;
    5447: romdata_int <= 'haee;
    5448: romdata_int <= 'h1c66;
    5449: romdata_int <= 'h414; // Line Descriptor
    5450: romdata_int <= 'h1800;
    5451: romdata_int <= 'hd2a;
    5452: romdata_int <= 'h1958;
    5453: romdata_int <= 'h414; // Line Descriptor
    5454: romdata_int <= 'h1a00;
    5455: romdata_int <= 'h1262;
    5456: romdata_int <= 'h12c1;
    5457: romdata_int <= 'h414; // Line Descriptor
    5458: romdata_int <= 'h1c00;
    5459: romdata_int <= 'h16b2;
    5460: romdata_int <= 'h79;
    5461: romdata_int <= 'h414; // Line Descriptor
    5462: romdata_int <= 'h1e00;
    5463: romdata_int <= 'h18e7;
    5464: romdata_int <= 'h231;
    5465: romdata_int <= 'h414; // Line Descriptor
    5466: romdata_int <= 'h2000;
    5467: romdata_int <= 'h1ea0;
    5468: romdata_int <= 'h6d0;
    5469: romdata_int <= 'h414; // Line Descriptor
    5470: romdata_int <= 'h2200;
    5471: romdata_int <= 'h1a30;
    5472: romdata_int <= 'h229b;
    5473: romdata_int <= 'h414; // Line Descriptor
    5474: romdata_int <= 'h2400;
    5475: romdata_int <= 'h4be;
    5476: romdata_int <= 'h2535;
    5477: romdata_int <= 'h414; // Line Descriptor
    5478: romdata_int <= 'h2600;
    5479: romdata_int <= 'h1cbd;
    5480: romdata_int <= 'h10c5;
    5481: romdata_int <= 'h414; // Line Descriptor
    5482: romdata_int <= 'h0;
    5483: romdata_int <= 'h209f;
    5484: romdata_int <= 'hd32;
    5485: romdata_int <= 'h414; // Line Descriptor
    5486: romdata_int <= 'h200;
    5487: romdata_int <= 'h1a1c;
    5488: romdata_int <= 'h125f;
    5489: romdata_int <= 'h414; // Line Descriptor
    5490: romdata_int <= 'h400;
    5491: romdata_int <= 'h142a;
    5492: romdata_int <= 'h1cc9;
    5493: romdata_int <= 'h414; // Line Descriptor
    5494: romdata_int <= 'h600;
    5495: romdata_int <= 'h519;
    5496: romdata_int <= 'h250;
    5497: romdata_int <= 'h414; // Line Descriptor
    5498: romdata_int <= 'h800;
    5499: romdata_int <= 'hb2c;
    5500: romdata_int <= 'h81a;
    5501: romdata_int <= 'h414; // Line Descriptor
    5502: romdata_int <= 'ha00;
    5503: romdata_int <= 'h1706;
    5504: romdata_int <= 'h721;
    5505: romdata_int <= 'h414; // Line Descriptor
    5506: romdata_int <= 'hc00;
    5507: romdata_int <= 'h1808;
    5508: romdata_int <= 'h1865;
    5509: romdata_int <= 'h414; // Line Descriptor
    5510: romdata_int <= 'he00;
    5511: romdata_int <= 'h1e5d;
    5512: romdata_int <= 'h1e7b;
    5513: romdata_int <= 'h414; // Line Descriptor
    5514: romdata_int <= 'h1000;
    5515: romdata_int <= 'h2218;
    5516: romdata_int <= 'h1640;
    5517: romdata_int <= 'h414; // Line Descriptor
    5518: romdata_int <= 'h1200;
    5519: romdata_int <= 'hc80;
    5520: romdata_int <= 'h14ab;
    5521: romdata_int <= 'h414; // Line Descriptor
    5522: romdata_int <= 'h1400;
    5523: romdata_int <= 'h123e;
    5524: romdata_int <= 'h25;
    5525: romdata_int <= 'h414; // Line Descriptor
    5526: romdata_int <= 'h1600;
    5527: romdata_int <= 'h893;
    5528: romdata_int <= 'h1061;
    5529: romdata_int <= 'h414; // Line Descriptor
    5530: romdata_int <= 'h1800;
    5531: romdata_int <= 'h1146;
    5532: romdata_int <= 'h2690;
    5533: romdata_int <= 'h414; // Line Descriptor
    5534: romdata_int <= 'h1a00;
    5535: romdata_int <= 'h670;
    5536: romdata_int <= 'h20b4;
    5537: romdata_int <= 'h414; // Line Descriptor
    5538: romdata_int <= 'h1c00;
    5539: romdata_int <= 'he2b;
    5540: romdata_int <= 'h1aba;
    5541: romdata_int <= 'h414; // Line Descriptor
    5542: romdata_int <= 'h1e00;
    5543: romdata_int <= 'h1c44;
    5544: romdata_int <= 'h4eb;
    5545: romdata_int <= 'h414; // Line Descriptor
    5546: romdata_int <= 'h2000;
    5547: romdata_int <= 'h24ea;
    5548: romdata_int <= 'ha72;
    5549: romdata_int <= 'h414; // Line Descriptor
    5550: romdata_int <= 'h2200;
    5551: romdata_int <= 'hee;
    5552: romdata_int <= 'h22c3;
    5553: romdata_int <= 'h414; // Line Descriptor
    5554: romdata_int <= 'h2400;
    5555: romdata_int <= 'h265c;
    5556: romdata_int <= 'h24ca;
    5557: romdata_int <= 'h414; // Line Descriptor
    5558: romdata_int <= 'h2600;
    5559: romdata_int <= 'h333;
    5560: romdata_int <= 'heb0;
    5561: romdata_int <= 'h414; // Line Descriptor
    5562: romdata_int <= 'h0;
    5563: romdata_int <= 'h106b;
    5564: romdata_int <= 'hcfd;
    5565: romdata_int <= 'h414; // Line Descriptor
    5566: romdata_int <= 'h200;
    5567: romdata_int <= 'hc41;
    5568: romdata_int <= 'ha07;
    5569: romdata_int <= 'h414; // Line Descriptor
    5570: romdata_int <= 'h400;
    5571: romdata_int <= 'h2673;
    5572: romdata_int <= 'h162b;
    5573: romdata_int <= 'h414; // Line Descriptor
    5574: romdata_int <= 'h600;
    5575: romdata_int <= 'h6ad;
    5576: romdata_int <= 'h235;
    5577: romdata_int <= 'h414; // Line Descriptor
    5578: romdata_int <= 'h800;
    5579: romdata_int <= 'h1d15;
    5580: romdata_int <= 'hf4c;
    5581: romdata_int <= 'h414; // Line Descriptor
    5582: romdata_int <= 'ha00;
    5583: romdata_int <= 'h2323;
    5584: romdata_int <= 'h2610;
    5585: romdata_int <= 'h414; // Line Descriptor
    5586: romdata_int <= 'hc00;
    5587: romdata_int <= 'h323;
    5588: romdata_int <= 'h18f6;
    5589: romdata_int <= 'h414; // Line Descriptor
    5590: romdata_int <= 'he00;
    5591: romdata_int <= 'h213d;
    5592: romdata_int <= 'h20ed;
    5593: romdata_int <= 'h414; // Line Descriptor
    5594: romdata_int <= 'h1000;
    5595: romdata_int <= 'h14c4;
    5596: romdata_int <= 'h2414;
    5597: romdata_int <= 'h414; // Line Descriptor
    5598: romdata_int <= 'h1200;
    5599: romdata_int <= 'h160a;
    5600: romdata_int <= 'h1c9a;
    5601: romdata_int <= 'h414; // Line Descriptor
    5602: romdata_int <= 'h1400;
    5603: romdata_int <= 'he32;
    5604: romdata_int <= 'h10f6;
    5605: romdata_int <= 'h414; // Line Descriptor
    5606: romdata_int <= 'h1600;
    5607: romdata_int <= 'h8b3;
    5608: romdata_int <= 'h1e3d;
    5609: romdata_int <= 'h414; // Line Descriptor
    5610: romdata_int <= 'h1800;
    5611: romdata_int <= 'h55d;
    5612: romdata_int <= 'h128f;
    5613: romdata_int <= 'h414; // Line Descriptor
    5614: romdata_int <= 'h1a00;
    5615: romdata_int <= 'h1850;
    5616: romdata_int <= 'h1a32;
    5617: romdata_int <= 'h414; // Line Descriptor
    5618: romdata_int <= 'h1c00;
    5619: romdata_int <= 'h1a2f;
    5620: romdata_int <= 'h8f8;
    5621: romdata_int <= 'h414; // Line Descriptor
    5622: romdata_int <= 'h1e00;
    5623: romdata_int <= 'h1ee3;
    5624: romdata_int <= 'h14dc;
    5625: romdata_int <= 'h414; // Line Descriptor
    5626: romdata_int <= 'h2000;
    5627: romdata_int <= 'haf6;
    5628: romdata_int <= 'h4f2;
    5629: romdata_int <= 'h414; // Line Descriptor
    5630: romdata_int <= 'h2200;
    5631: romdata_int <= 'h2520;
    5632: romdata_int <= 'h1e;
    5633: romdata_int <= 'h414; // Line Descriptor
    5634: romdata_int <= 'h2400;
    5635: romdata_int <= 'h1345;
    5636: romdata_int <= 'h2278;
    5637: romdata_int <= 'h414; // Line Descriptor
    5638: romdata_int <= 'h2600;
    5639: romdata_int <= 'h3f;
    5640: romdata_int <= 'h6f5;
    5641: romdata_int <= 'h414; // Line Descriptor
    5642: romdata_int <= 'h0;
    5643: romdata_int <= 'h12a8;
    5644: romdata_int <= 'h1697;
    5645: romdata_int <= 'h414; // Line Descriptor
    5646: romdata_int <= 'h200;
    5647: romdata_int <= 'h22b1;
    5648: romdata_int <= 'h8a1;
    5649: romdata_int <= 'h414; // Line Descriptor
    5650: romdata_int <= 'h400;
    5651: romdata_int <= 'h1097;
    5652: romdata_int <= 'h61d;
    5653: romdata_int <= 'h414; // Line Descriptor
    5654: romdata_int <= 'h600;
    5655: romdata_int <= 'h24a2;
    5656: romdata_int <= 'h16;
    5657: romdata_int <= 'h414; // Line Descriptor
    5658: romdata_int <= 'h800;
    5659: romdata_int <= 'hd37;
    5660: romdata_int <= 'h1f4c;
    5661: romdata_int <= 'h414; // Line Descriptor
    5662: romdata_int <= 'ha00;
    5663: romdata_int <= 'h1ef4;
    5664: romdata_int <= 'h1c36;
    5665: romdata_int <= 'h414; // Line Descriptor
    5666: romdata_int <= 'hc00;
    5667: romdata_int <= 'h24a;
    5668: romdata_int <= 'hf56;
    5669: romdata_int <= 'h414; // Line Descriptor
    5670: romdata_int <= 'he00;
    5671: romdata_int <= 'h1add;
    5672: romdata_int <= 'h1860;
    5673: romdata_int <= 'h414; // Line Descriptor
    5674: romdata_int <= 'h1000;
    5675: romdata_int <= 'he69;
    5676: romdata_int <= 'h1252;
    5677: romdata_int <= 'h414; // Line Descriptor
    5678: romdata_int <= 'h1200;
    5679: romdata_int <= 'h2669;
    5680: romdata_int <= 'ha67;
    5681: romdata_int <= 'h414; // Line Descriptor
    5682: romdata_int <= 'h1400;
    5683: romdata_int <= 'h6c8;
    5684: romdata_int <= 'h113f;
    5685: romdata_int <= 'h414; // Line Descriptor
    5686: romdata_int <= 'h1600;
    5687: romdata_int <= 'h150;
    5688: romdata_int <= 'h4b5;
    5689: romdata_int <= 'h414; // Line Descriptor
    5690: romdata_int <= 'h1800;
    5691: romdata_int <= 'h1cb8;
    5692: romdata_int <= 'h2e2;
    5693: romdata_int <= 'h414; // Line Descriptor
    5694: romdata_int <= 'h1a00;
    5695: romdata_int <= 'h83a;
    5696: romdata_int <= 'h1560;
    5697: romdata_int <= 'h414; // Line Descriptor
    5698: romdata_int <= 'h1c00;
    5699: romdata_int <= 'ha62;
    5700: romdata_int <= 'h1ab4;
    5701: romdata_int <= 'h414; // Line Descriptor
    5702: romdata_int <= 'h1e00;
    5703: romdata_int <= 'h16d8;
    5704: romdata_int <= 'hc03;
    5705: romdata_int <= 'h414; // Line Descriptor
    5706: romdata_int <= 'h2000;
    5707: romdata_int <= 'h1494;
    5708: romdata_int <= 'h2059;
    5709: romdata_int <= 'h414; // Line Descriptor
    5710: romdata_int <= 'h2200;
    5711: romdata_int <= 'h18e8;
    5712: romdata_int <= 'h24a0;
    5713: romdata_int <= 'h414; // Line Descriptor
    5714: romdata_int <= 'h2400;
    5715: romdata_int <= 'h458;
    5716: romdata_int <= 'h22ee;
    5717: romdata_int <= 'h414; // Line Descriptor
    5718: romdata_int <= 'h2600;
    5719: romdata_int <= 'h211e;
    5720: romdata_int <= 'h2645;
    5721: romdata_int <= 'h414; // Line Descriptor
    5722: romdata_int <= 'h0;
    5723: romdata_int <= 'h1430;
    5724: romdata_int <= 'h1880;
    5725: romdata_int <= 'h414; // Line Descriptor
    5726: romdata_int <= 'h200;
    5727: romdata_int <= 'h467;
    5728: romdata_int <= 'h2749;
    5729: romdata_int <= 'h414; // Line Descriptor
    5730: romdata_int <= 'h400;
    5731: romdata_int <= 'h22e5;
    5732: romdata_int <= 'h14f3;
    5733: romdata_int <= 'h414; // Line Descriptor
    5734: romdata_int <= 'h600;
    5735: romdata_int <= 'h103d;
    5736: romdata_int <= 'h1b59;
    5737: romdata_int <= 'h414; // Line Descriptor
    5738: romdata_int <= 'h800;
    5739: romdata_int <= 'h26cf;
    5740: romdata_int <= 'h2233;
    5741: romdata_int <= 'h414; // Line Descriptor
    5742: romdata_int <= 'ha00;
    5743: romdata_int <= 'h2091;
    5744: romdata_int <= 'h476;
    5745: romdata_int <= 'h414; // Line Descriptor
    5746: romdata_int <= 'hc00;
    5747: romdata_int <= 'h1e13;
    5748: romdata_int <= 'hc3d;
    5749: romdata_int <= 'h414; // Line Descriptor
    5750: romdata_int <= 'he00;
    5751: romdata_int <= 'h1759;
    5752: romdata_int <= 'h10e3;
    5753: romdata_int <= 'h414; // Line Descriptor
    5754: romdata_int <= 'h1000;
    5755: romdata_int <= 'h24e6;
    5756: romdata_int <= 'h270;
    5757: romdata_int <= 'h414; // Line Descriptor
    5758: romdata_int <= 'h1200;
    5759: romdata_int <= 'hce;
    5760: romdata_int <= 'hd6;
    5761: romdata_int <= 'h414; // Line Descriptor
    5762: romdata_int <= 'h1400;
    5763: romdata_int <= 'hb23;
    5764: romdata_int <= 'h1c17;
    5765: romdata_int <= 'h414; // Line Descriptor
    5766: romdata_int <= 'h1600;
    5767: romdata_int <= 'h1c6b;
    5768: romdata_int <= 'h2515;
    5769: romdata_int <= 'h414; // Line Descriptor
    5770: romdata_int <= 'h1800;
    5771: romdata_int <= 'h1abd;
    5772: romdata_int <= 'h1711;
    5773: romdata_int <= 'h414; // Line Descriptor
    5774: romdata_int <= 'h1a00;
    5775: romdata_int <= 'hf1d;
    5776: romdata_int <= 'h1e4f;
    5777: romdata_int <= 'h414; // Line Descriptor
    5778: romdata_int <= 'h1c00;
    5779: romdata_int <= 'h646;
    5780: romdata_int <= 'ha10;
    5781: romdata_int <= 'h414; // Line Descriptor
    5782: romdata_int <= 'h1e00;
    5783: romdata_int <= 'h34a;
    5784: romdata_int <= 'h703;
    5785: romdata_int <= 'h414; // Line Descriptor
    5786: romdata_int <= 'h2000;
    5787: romdata_int <= 'h133e;
    5788: romdata_int <= 'h12e4;
    5789: romdata_int <= 'h414; // Line Descriptor
    5790: romdata_int <= 'h2200;
    5791: romdata_int <= 'hcf2;
    5792: romdata_int <= 'h202c;
    5793: romdata_int <= 'h414; // Line Descriptor
    5794: romdata_int <= 'h2400;
    5795: romdata_int <= 'h1962;
    5796: romdata_int <= 'h935;
    5797: romdata_int <= 'h414; // Line Descriptor
    5798: romdata_int <= 'h2600;
    5799: romdata_int <= 'h952;
    5800: romdata_int <= 'hf64;
    5801: romdata_int <= 'h414; // Line Descriptor
    5802: romdata_int <= 'h0;
    5803: romdata_int <= 'h253d;
    5804: romdata_int <= 'h1661;
    5805: romdata_int <= 'h414; // Line Descriptor
    5806: romdata_int <= 'h200;
    5807: romdata_int <= 'h229b;
    5808: romdata_int <= 'h15c;
    5809: romdata_int <= 'h414; // Line Descriptor
    5810: romdata_int <= 'h400;
    5811: romdata_int <= 'h1487;
    5812: romdata_int <= 'h561;
    5813: romdata_int <= 'h414; // Line Descriptor
    5814: romdata_int <= 'h600;
    5815: romdata_int <= 'h1a38;
    5816: romdata_int <= 'h8b4;
    5817: romdata_int <= 'h414; // Line Descriptor
    5818: romdata_int <= 'h800;
    5819: romdata_int <= 'h1cb8;
    5820: romdata_int <= 'h2220;
    5821: romdata_int <= 'h414; // Line Descriptor
    5822: romdata_int <= 'ha00;
    5823: romdata_int <= 'h1e43;
    5824: romdata_int <= 'h1405;
    5825: romdata_int <= 'h414; // Line Descriptor
    5826: romdata_int <= 'hc00;
    5827: romdata_int <= 'h12a6;
    5828: romdata_int <= 'h2150;
    5829: romdata_int <= 'h414; // Line Descriptor
    5830: romdata_int <= 'he00;
    5831: romdata_int <= 'ha7d;
    5832: romdata_int <= 'heaa;
    5833: romdata_int <= 'h414; // Line Descriptor
    5834: romdata_int <= 'h1000;
    5835: romdata_int <= 'h47b;
    5836: romdata_int <= 'hcf0;
    5837: romdata_int <= 'h414; // Line Descriptor
    5838: romdata_int <= 'h1200;
    5839: romdata_int <= 'h20d2;
    5840: romdata_int <= 'h1c0a;
    5841: romdata_int <= 'h414; // Line Descriptor
    5842: romdata_int <= 'h1400;
    5843: romdata_int <= 'h110b;
    5844: romdata_int <= 'h2718;
    5845: romdata_int <= 'h414; // Line Descriptor
    5846: romdata_int <= 'h1600;
    5847: romdata_int <= 'hf4b;
    5848: romdata_int <= 'h738;
    5849: romdata_int <= 'h414; // Line Descriptor
    5850: romdata_int <= 'h1800;
    5851: romdata_int <= 'h884;
    5852: romdata_int <= 'h1afd;
    5853: romdata_int <= 'h414; // Line Descriptor
    5854: romdata_int <= 'h1a00;
    5855: romdata_int <= 'h18d2;
    5856: romdata_int <= 'h10fe;
    5857: romdata_int <= 'h414; // Line Descriptor
    5858: romdata_int <= 'h1c00;
    5859: romdata_int <= 'h6ad;
    5860: romdata_int <= 'h12c2;
    5861: romdata_int <= 'h414; // Line Descriptor
    5862: romdata_int <= 'h1e00;
    5863: romdata_int <= 'hd09;
    5864: romdata_int <= 'h2417;
    5865: romdata_int <= 'h414; // Line Descriptor
    5866: romdata_int <= 'h2000;
    5867: romdata_int <= 'hd8;
    5868: romdata_int <= 'h332;
    5869: romdata_int <= 'h414; // Line Descriptor
    5870: romdata_int <= 'h2200;
    5871: romdata_int <= 'h2c6;
    5872: romdata_int <= 'ha38;
    5873: romdata_int <= 'h414; // Line Descriptor
    5874: romdata_int <= 'h2400;
    5875: romdata_int <= 'h271c;
    5876: romdata_int <= 'h1e3b;
    5877: romdata_int <= 'h414; // Line Descriptor
    5878: romdata_int <= 'h2600;
    5879: romdata_int <= 'h1745;
    5880: romdata_int <= 'h1827;
    5881: romdata_int <= 'h414; // Line Descriptor
    5882: romdata_int <= 'h0;
    5883: romdata_int <= 'h1cc4;
    5884: romdata_int <= 'h248a;
    5885: romdata_int <= 'h414; // Line Descriptor
    5886: romdata_int <= 'h200;
    5887: romdata_int <= 'h24a1;
    5888: romdata_int <= 'hf49;
    5889: romdata_int <= 'h414; // Line Descriptor
    5890: romdata_int <= 'h400;
    5891: romdata_int <= 'h1637;
    5892: romdata_int <= 'h2149;
    5893: romdata_int <= 'h414; // Line Descriptor
    5894: romdata_int <= 'h600;
    5895: romdata_int <= 'h2248;
    5896: romdata_int <= 'hd37;
    5897: romdata_int <= 'h414; // Line Descriptor
    5898: romdata_int <= 'h800;
    5899: romdata_int <= 'hc48;
    5900: romdata_int <= 'hac2;
    5901: romdata_int <= 'h414; // Line Descriptor
    5902: romdata_int <= 'ha00;
    5903: romdata_int <= 'hec3;
    5904: romdata_int <= 'h6ca;
    5905: romdata_int <= 'h414; // Line Descriptor
    5906: romdata_int <= 'hc00;
    5907: romdata_int <= 'h2755;
    5908: romdata_int <= 'h1a8f;
    5909: romdata_int <= 'h414; // Line Descriptor
    5910: romdata_int <= 'he00;
    5911: romdata_int <= 'h1a56;
    5912: romdata_int <= 'h1f18;
    5913: romdata_int <= 'h414; // Line Descriptor
    5914: romdata_int <= 'h1000;
    5915: romdata_int <= 'h504;
    5916: romdata_int <= 'h12d5;
    5917: romdata_int <= 'h414; // Line Descriptor
    5918: romdata_int <= 'h1200;
    5919: romdata_int <= 'h897;
    5920: romdata_int <= 'h4ec;
    5921: romdata_int <= 'h414; // Line Descriptor
    5922: romdata_int <= 'h1400;
    5923: romdata_int <= 'hb10;
    5924: romdata_int <= 'h193e;
    5925: romdata_int <= 'h414; // Line Descriptor
    5926: romdata_int <= 'h1600;
    5927: romdata_int <= 'h1412;
    5928: romdata_int <= 'h105b;
    5929: romdata_int <= 'h414; // Line Descriptor
    5930: romdata_int <= 'h1800;
    5931: romdata_int <= 'h1eea;
    5932: romdata_int <= 'h50;
    5933: romdata_int <= 'h414; // Line Descriptor
    5934: romdata_int <= 'h1a00;
    5935: romdata_int <= 'h22;
    5936: romdata_int <= 'h1c67;
    5937: romdata_int <= 'h414; // Line Descriptor
    5938: romdata_int <= 'h1c00;
    5939: romdata_int <= 'h25a;
    5940: romdata_int <= 'h154e;
    5941: romdata_int <= 'h414; // Line Descriptor
    5942: romdata_int <= 'h1e00;
    5943: romdata_int <= 'h1285;
    5944: romdata_int <= 'h2244;
    5945: romdata_int <= 'h414; // Line Descriptor
    5946: romdata_int <= 'h2000;
    5947: romdata_int <= 'h67b;
    5948: romdata_int <= 'h254;
    5949: romdata_int <= 'h414; // Line Descriptor
    5950: romdata_int <= 'h2200;
    5951: romdata_int <= 'h192a;
    5952: romdata_int <= 'h1702;
    5953: romdata_int <= 'h414; // Line Descriptor
    5954: romdata_int <= 'h2400;
    5955: romdata_int <= 'h111e;
    5956: romdata_int <= 'h8d6;
    5957: romdata_int <= 'h514; // Line Descriptor
    5958: romdata_int <= 'h2600;
    5959: romdata_int <= 'h2054;
    5960: romdata_int <= 'h2648;
    5961: romdata_int <= 'h612; // Line Descriptor
    5962: romdata_int <= 'h0;
    5963: romdata_int <= 'h1b37;
    5964: romdata_int <= 'he8e;
    5965: romdata_int <= 'h4a1;
    5966: romdata_int <= 'h612; // Line Descriptor
    5967: romdata_int <= 'h200;
    5968: romdata_int <= 'h122;
    5969: romdata_int <= 'h16ae;
    5970: romdata_int <= 'hf0b;
    5971: romdata_int <= 'h612; // Line Descriptor
    5972: romdata_int <= 'h400;
    5973: romdata_int <= 'h1e89;
    5974: romdata_int <= 'hc2e;
    5975: romdata_int <= 'h1204;
    5976: romdata_int <= 'h612; // Line Descriptor
    5977: romdata_int <= 'h600;
    5978: romdata_int <= 'h35c;
    5979: romdata_int <= 'h1ce1;
    5980: romdata_int <= 'h22ec;
    5981: romdata_int <= 'h612; // Line Descriptor
    5982: romdata_int <= 'h800;
    5983: romdata_int <= 'h163a;
    5984: romdata_int <= 'h20a1;
    5985: romdata_int <= 'h939;
    5986: romdata_int <= 'h612; // Line Descriptor
    5987: romdata_int <= 'ha00;
    5988: romdata_int <= 'hc60;
    5989: romdata_int <= 'h879;
    5990: romdata_int <= 'h6b8;
    5991: romdata_int <= 'h612; // Line Descriptor
    5992: romdata_int <= 'hc00;
    5993: romdata_int <= 'h18b9;
    5994: romdata_int <= 'h113b;
    5995: romdata_int <= 'h1c7c;
    5996: romdata_int <= 'h612; // Line Descriptor
    5997: romdata_int <= 'he00;
    5998: romdata_int <= 'he79;
    5999: romdata_int <= 'h181e;
    6000: romdata_int <= 'h2bc;
    6001: romdata_int <= 'h612; // Line Descriptor
    6002: romdata_int <= 'h1000;
    6003: romdata_int <= 'ha91;
    6004: romdata_int <= 'h40d;
    6005: romdata_int <= 'hd28;
    6006: romdata_int <= 'h612; // Line Descriptor
    6007: romdata_int <= 'h1200;
    6008: romdata_int <= 'h2055;
    6009: romdata_int <= 'h1261;
    6010: romdata_int <= 'h18d5;
    6011: romdata_int <= 'h612; // Line Descriptor
    6012: romdata_int <= 'h1400;
    6013: romdata_int <= 'h1ce6;
    6014: romdata_int <= 'h2334;
    6015: romdata_int <= 'h14ae;
    6016: romdata_int <= 'h612; // Line Descriptor
    6017: romdata_int <= 'h1600;
    6018: romdata_int <= 'h10f3;
    6019: romdata_int <= 'haa4;
    6020: romdata_int <= 'h12c;
    6021: romdata_int <= 'h612; // Line Descriptor
    6022: romdata_int <= 'h1800;
    6023: romdata_int <= 'h643;
    6024: romdata_int <= 'h328;
    6025: romdata_int <= 'h16b0;
    6026: romdata_int <= 'h612; // Line Descriptor
    6027: romdata_int <= 'h1a00;
    6028: romdata_int <= 'h224e;
    6029: romdata_int <= 'hc4;
    6030: romdata_int <= 'h1f50;
    6031: romdata_int <= 'h612; // Line Descriptor
    6032: romdata_int <= 'h1c00;
    6033: romdata_int <= 'h852;
    6034: romdata_int <= 'h143b;
    6035: romdata_int <= 'h212b;
    6036: romdata_int <= 'h612; // Line Descriptor
    6037: romdata_int <= 'h1e00;
    6038: romdata_int <= 'h12d5;
    6039: romdata_int <= 'h1a62;
    6040: romdata_int <= 'h1af2;
    6041: romdata_int <= 'h612; // Line Descriptor
    6042: romdata_int <= 'h2000;
    6043: romdata_int <= 'h44a;
    6044: romdata_int <= 'h677;
    6045: romdata_int <= 'hae7;
    6046: romdata_int <= 'h612; // Line Descriptor
    6047: romdata_int <= 'h2200;
    6048: romdata_int <= 'h1483;
    6049: romdata_int <= 'h1f18;
    6050: romdata_int <= 'h100e;
    6051: romdata_int <= 'h412; // Line Descriptor
    6052: romdata_int <= 'h0;
    6053: romdata_int <= 'h2153;
    6054: romdata_int <= 'hb2c;
    6055: romdata_int <= 'h412; // Line Descriptor
    6056: romdata_int <= 'h200;
    6057: romdata_int <= 'hca6;
    6058: romdata_int <= 'h1cf2;
    6059: romdata_int <= 'h412; // Line Descriptor
    6060: romdata_int <= 'h400;
    6061: romdata_int <= 'h6bd;
    6062: romdata_int <= 'h1a5c;
    6063: romdata_int <= 'h412; // Line Descriptor
    6064: romdata_int <= 'h600;
    6065: romdata_int <= 'h1d01;
    6066: romdata_int <= 'hd34;
    6067: romdata_int <= 'h412; // Line Descriptor
    6068: romdata_int <= 'h800;
    6069: romdata_int <= 'h84b;
    6070: romdata_int <= 'h1ed9;
    6071: romdata_int <= 'h412; // Line Descriptor
    6072: romdata_int <= 'ha00;
    6073: romdata_int <= 'h1206;
    6074: romdata_int <= 'h65f;
    6075: romdata_int <= 'h412; // Line Descriptor
    6076: romdata_int <= 'hc00;
    6077: romdata_int <= 'hf2d;
    6078: romdata_int <= 'h89f;
    6079: romdata_int <= 'h412; // Line Descriptor
    6080: romdata_int <= 'he00;
    6081: romdata_int <= 'h234f;
    6082: romdata_int <= 'h2225;
    6083: romdata_int <= 'h412; // Line Descriptor
    6084: romdata_int <= 'h1000;
    6085: romdata_int <= 'h138;
    6086: romdata_int <= 'h108f;
    6087: romdata_int <= 'h412; // Line Descriptor
    6088: romdata_int <= 'h1200;
    6089: romdata_int <= 'h475;
    6090: romdata_int <= 'h1241;
    6091: romdata_int <= 'h412; // Line Descriptor
    6092: romdata_int <= 'h1400;
    6093: romdata_int <= 'h1e33;
    6094: romdata_int <= 'hf11;
    6095: romdata_int <= 'h412; // Line Descriptor
    6096: romdata_int <= 'h1600;
    6097: romdata_int <= 'h1b4a;
    6098: romdata_int <= 'h167d;
    6099: romdata_int <= 'h412; // Line Descriptor
    6100: romdata_int <= 'h1800;
    6101: romdata_int <= 'h104f;
    6102: romdata_int <= 'h305;
    6103: romdata_int <= 'h412; // Line Descriptor
    6104: romdata_int <= 'h1a00;
    6105: romdata_int <= 'h348;
    6106: romdata_int <= 'h181a;
    6107: romdata_int <= 'h412; // Line Descriptor
    6108: romdata_int <= 'h1c00;
    6109: romdata_int <= 'haee;
    6110: romdata_int <= 'h1466;
    6111: romdata_int <= 'h412; // Line Descriptor
    6112: romdata_int <= 'h1e00;
    6113: romdata_int <= 'h152a;
    6114: romdata_int <= 'h2158;
    6115: romdata_int <= 'h412; // Line Descriptor
    6116: romdata_int <= 'h2000;
    6117: romdata_int <= 'h1662;
    6118: romdata_int <= 'h4c1;
    6119: romdata_int <= 'h412; // Line Descriptor
    6120: romdata_int <= 'h2200;
    6121: romdata_int <= 'h18b2;
    6122: romdata_int <= 'h79;
    6123: romdata_int <= 'h412; // Line Descriptor
    6124: romdata_int <= 'h0;
    6125: romdata_int <= 'hee7;
    6126: romdata_int <= 'h431;
    6127: romdata_int <= 'h412; // Line Descriptor
    6128: romdata_int <= 'h200;
    6129: romdata_int <= 'h20a0;
    6130: romdata_int <= 'hd0;
    6131: romdata_int <= 'h412; // Line Descriptor
    6132: romdata_int <= 'h400;
    6133: romdata_int <= 'h1430;
    6134: romdata_int <= 'h169b;
    6135: romdata_int <= 'h412; // Line Descriptor
    6136: romdata_int <= 'h600;
    6137: romdata_int <= 'h6be;
    6138: romdata_int <= 'h2335;
    6139: romdata_int <= 'h412; // Line Descriptor
    6140: romdata_int <= 'h800;
    6141: romdata_int <= 'h4bd;
    6142: romdata_int <= 'hcc5;
    6143: romdata_int <= 'h412; // Line Descriptor
    6144: romdata_int <= 'ha00;
    6145: romdata_int <= 'h1c9f;
    6146: romdata_int <= 'hf32;
    6147: romdata_int <= 'h412; // Line Descriptor
    6148: romdata_int <= 'hc00;
    6149: romdata_int <= 'h181c;
    6150: romdata_int <= 'h125f;
    6151: romdata_int <= 'h412; // Line Descriptor
    6152: romdata_int <= 'he00;
    6153: romdata_int <= 'h122a;
    6154: romdata_int <= 'h1ac9;
    6155: romdata_int <= 'h412; // Line Descriptor
    6156: romdata_int <= 'h1000;
    6157: romdata_int <= 'h319;
    6158: romdata_int <= 'h250;
    6159: romdata_int <= 'h412; // Line Descriptor
    6160: romdata_int <= 'h1200;
    6161: romdata_int <= 'h1b38;
    6162: romdata_int <= 'h821;
    6163: romdata_int <= 'h412; // Line Descriptor
    6164: romdata_int <= 'h1400;
    6165: romdata_int <= 'hb2c;
    6166: romdata_int <= 'ha1a;
    6167: romdata_int <= 'h412; // Line Descriptor
    6168: romdata_int <= 'h1600;
    6169: romdata_int <= 'h1106;
    6170: romdata_int <= 'h1121;
    6171: romdata_int <= 'h412; // Line Descriptor
    6172: romdata_int <= 'h1800;
    6173: romdata_int <= 'h1608;
    6174: romdata_int <= 'h1c65;
    6175: romdata_int <= 'h412; // Line Descriptor
    6176: romdata_int <= 'h1a00;
    6177: romdata_int <= 'h1e5d;
    6178: romdata_int <= 'h1e7b;
    6179: romdata_int <= 'h412; // Line Descriptor
    6180: romdata_int <= 'h1c00;
    6181: romdata_int <= 'h2218;
    6182: romdata_int <= 'h1840;
    6183: romdata_int <= 'h412; // Line Descriptor
    6184: romdata_int <= 'h1e00;
    6185: romdata_int <= 'h880;
    6186: romdata_int <= 'h14ab;
    6187: romdata_int <= 'h412; // Line Descriptor
    6188: romdata_int <= 'h2000;
    6189: romdata_int <= 'hc3e;
    6190: romdata_int <= 'h625;
    6191: romdata_int <= 'h412; // Line Descriptor
    6192: romdata_int <= 'h2200;
    6193: romdata_int <= 'h7e;
    6194: romdata_int <= 'h213f;
    6195: romdata_int <= 'h412; // Line Descriptor
    6196: romdata_int <= 'h0;
    6197: romdata_int <= 'h1546;
    6198: romdata_int <= 'h2290;
    6199: romdata_int <= 'h412; // Line Descriptor
    6200: romdata_int <= 'h200;
    6201: romdata_int <= 'h102b;
    6202: romdata_int <= 'h16ba;
    6203: romdata_int <= 'h412; // Line Descriptor
    6204: romdata_int <= 'h400;
    6205: romdata_int <= 'he44;
    6206: romdata_int <= 'h2eb;
    6207: romdata_int <= 'h412; // Line Descriptor
    6208: romdata_int <= 'h600;
    6209: romdata_int <= 'h1aea;
    6210: romdata_int <= 'h72;
    6211: romdata_int <= 'h412; // Line Descriptor
    6212: romdata_int <= 'h800;
    6213: romdata_int <= 'h4ee;
    6214: romdata_int <= 'hec3;
    6215: romdata_int <= 'h412; // Line Descriptor
    6216: romdata_int <= 'ha00;
    6217: romdata_int <= 'hb33;
    6218: romdata_int <= 'h20b0;
    6219: romdata_int <= 'h412; // Line Descriptor
    6220: romdata_int <= 'hc00;
    6221: romdata_int <= 'h126b;
    6222: romdata_int <= 'hcfd;
    6223: romdata_int <= 'h412; // Line Descriptor
    6224: romdata_int <= 'he00;
    6225: romdata_int <= 'h841;
    6226: romdata_int <= 'ha07;
    6227: romdata_int <= 'h412; // Line Descriptor
    6228: romdata_int <= 'h1000;
    6229: romdata_int <= 'h2ad;
    6230: romdata_int <= 'h435;
    6231: romdata_int <= 'h412; // Line Descriptor
    6232: romdata_int <= 'h1200;
    6233: romdata_int <= 'h1ead;
    6234: romdata_int <= 'h103c;
    6235: romdata_int <= 'h412; // Line Descriptor
    6236: romdata_int <= 'h1400;
    6237: romdata_int <= 'h123;
    6238: romdata_int <= 'h18f6;
    6239: romdata_int <= 'h412; // Line Descriptor
    6240: romdata_int <= 'h1600;
    6241: romdata_int <= 'h213d;
    6242: romdata_int <= 'h1ced;
    6243: romdata_int <= 'h412; // Line Descriptor
    6244: romdata_int <= 'h1800;
    6245: romdata_int <= 'h18c4;
    6246: romdata_int <= 'h1e14;
    6247: romdata_int <= 'h412; // Line Descriptor
    6248: romdata_int <= 'h1a00;
    6249: romdata_int <= 'h160a;
    6250: romdata_int <= 'h149a;
    6251: romdata_int <= 'h412; // Line Descriptor
    6252: romdata_int <= 'h1c00;
    6253: romdata_int <= 'hc32;
    6254: romdata_int <= 'h8f6;
    6255: romdata_int <= 'h412; // Line Descriptor
    6256: romdata_int <= 'h1e00;
    6257: romdata_int <= 'h6b3;
    6258: romdata_int <= 'h1a3d;
    6259: romdata_int <= 'h412; // Line Descriptor
    6260: romdata_int <= 'h2000;
    6261: romdata_int <= 'h1d5d;
    6262: romdata_int <= 'h128f;
    6263: romdata_int <= 'h412; // Line Descriptor
    6264: romdata_int <= 'h2200;
    6265: romdata_int <= 'h2250;
    6266: romdata_int <= 'h632;
    6267: romdata_int <= 'h412; // Line Descriptor
    6268: romdata_int <= 'h0;
    6269: romdata_int <= 'h122f;
    6270: romdata_int <= 'h16f8;
    6271: romdata_int <= 'h412; // Line Descriptor
    6272: romdata_int <= 'h200;
    6273: romdata_int <= 'h16e3;
    6274: romdata_int <= 'h14dc;
    6275: romdata_int <= 'h412; // Line Descriptor
    6276: romdata_int <= 'h400;
    6277: romdata_int <= 'haf6;
    6278: romdata_int <= 'haf2;
    6279: romdata_int <= 'h412; // Line Descriptor
    6280: romdata_int <= 'h600;
    6281: romdata_int <= 'h1d20;
    6282: romdata_int <= 'h21e;
    6283: romdata_int <= 'h412; // Line Descriptor
    6284: romdata_int <= 'h800;
    6285: romdata_int <= 'h183f;
    6286: romdata_int <= 'h20f5;
    6287: romdata_int <= 'h412; // Line Descriptor
    6288: romdata_int <= 'ha00;
    6289: romdata_int <= 'h20b1;
    6290: romdata_int <= 'h8a1;
    6291: romdata_int <= 'h412; // Line Descriptor
    6292: romdata_int <= 'hc00;
    6293: romdata_int <= 'hc97;
    6294: romdata_int <= 'h61d;
    6295: romdata_int <= 'h412; // Line Descriptor
    6296: romdata_int <= 'he00;
    6297: romdata_int <= 'h63c;
    6298: romdata_int <= 'h4e5;
    6299: romdata_int <= 'h412; // Line Descriptor
    6300: romdata_int <= 'h1000;
    6301: romdata_int <= 'h881;
    6302: romdata_int <= 'h134d;
    6303: romdata_int <= 'h412; // Line Descriptor
    6304: romdata_int <= 'h1200;
    6305: romdata_int <= 'hf37;
    6306: romdata_int <= 'h1d4c;
    6307: romdata_int <= 'h412; // Line Descriptor
    6308: romdata_int <= 'h1400;
    6309: romdata_int <= 'h4f3;
    6310: romdata_int <= 'h1a57;
    6311: romdata_int <= 'h412; // Line Descriptor
    6312: romdata_int <= 'h1600;
    6313: romdata_int <= 'h1ef4;
    6314: romdata_int <= 'h1836;
    6315: romdata_int <= 'h412; // Line Descriptor
    6316: romdata_int <= 'h1800;
    6317: romdata_int <= 'h4a;
    6318: romdata_int <= 'hf56;
    6319: romdata_int <= 'h412; // Line Descriptor
    6320: romdata_int <= 'h1a00;
    6321: romdata_int <= 'h1b29;
    6322: romdata_int <= 'h1edc;
    6323: romdata_int <= 'h412; // Line Descriptor
    6324: romdata_int <= 'h1c00;
    6325: romdata_int <= 'h2269;
    6326: romdata_int <= 'h67;
    6327: romdata_int <= 'h412; // Line Descriptor
    6328: romdata_int <= 'h1e00;
    6329: romdata_int <= 'h2c8;
    6330: romdata_int <= 'hd3f;
    6331: romdata_int <= 'h412; // Line Descriptor
    6332: romdata_int <= 'h2000;
    6333: romdata_int <= 'h1150;
    6334: romdata_int <= 'h10b5;
    6335: romdata_int <= 'h412; // Line Descriptor
    6336: romdata_int <= 'h2200;
    6337: romdata_int <= 'h14b8;
    6338: romdata_int <= 'h22e2;
    6339: romdata_int <= 'h412; // Line Descriptor
    6340: romdata_int <= 'h0;
    6341: romdata_int <= 'h862;
    6342: romdata_int <= 'h8b4;
    6343: romdata_int <= 'h412; // Line Descriptor
    6344: romdata_int <= 'h200;
    6345: romdata_int <= 'he77;
    6346: romdata_int <= 'h8;
    6347: romdata_int <= 'h412; // Line Descriptor
    6348: romdata_int <= 'h400;
    6349: romdata_int <= 'ha58;
    6350: romdata_int <= 'heee;
    6351: romdata_int <= 'h412; // Line Descriptor
    6352: romdata_int <= 'h600;
    6353: romdata_int <= 'hd1e;
    6354: romdata_int <= 'h1445;
    6355: romdata_int <= 'h412; // Line Descriptor
    6356: romdata_int <= 'h800;
    6357: romdata_int <= 'h267;
    6358: romdata_int <= 'h2349;
    6359: romdata_int <= 'h412; // Line Descriptor
    6360: romdata_int <= 'ha00;
    6361: romdata_int <= 'h1d0b;
    6362: romdata_int <= 'hc96;
    6363: romdata_int <= 'h412; // Line Descriptor
    6364: romdata_int <= 'hc00;
    6365: romdata_int <= 'h2251;
    6366: romdata_int <= 'h18ba;
    6367: romdata_int <= 'h412; // Line Descriptor
    6368: romdata_int <= 'he00;
    6369: romdata_int <= 'hed;
    6370: romdata_int <= 'h1226;
    6371: romdata_int <= 'h412; // Line Descriptor
    6372: romdata_int <= 'h1000;
    6373: romdata_int <= 'h20e6;
    6374: romdata_int <= 'h470;
    6375: romdata_int <= 'h412; // Line Descriptor
    6376: romdata_int <= 'h1200;
    6377: romdata_int <= 'h1e74;
    6378: romdata_int <= 'h1c29;
    6379: romdata_int <= 'h412; // Line Descriptor
    6380: romdata_int <= 'h1400;
    6381: romdata_int <= 'h4ce;
    6382: romdata_int <= 'h2d6;
    6383: romdata_int <= 'h412; // Line Descriptor
    6384: romdata_int <= 'h1600;
    6385: romdata_int <= 'h171c;
    6386: romdata_int <= 'h1a33;
    6387: romdata_int <= 'h412; // Line Descriptor
    6388: romdata_int <= 'h1800;
    6389: romdata_int <= 'h1155;
    6390: romdata_int <= 'h16b8;
    6391: romdata_int <= 'h412; // Line Descriptor
    6392: romdata_int <= 'h1a00;
    6393: romdata_int <= 'h1a6b;
    6394: romdata_int <= 'h2115;
    6395: romdata_int <= 'h412; // Line Descriptor
    6396: romdata_int <= 'h1c00;
    6397: romdata_int <= 'h151d;
    6398: romdata_int <= 'h1e4f;
    6399: romdata_int <= 'h412; // Line Descriptor
    6400: romdata_int <= 'h1e00;
    6401: romdata_int <= 'h646;
    6402: romdata_int <= 'ha10;
    6403: romdata_int <= 'h412; // Line Descriptor
    6404: romdata_int <= 'h2000;
    6405: romdata_int <= 'h134a;
    6406: romdata_int <= 'h703;
    6407: romdata_int <= 'h412; // Line Descriptor
    6408: romdata_int <= 'h2200;
    6409: romdata_int <= 'h18fc;
    6410: romdata_int <= 'h1162;
    6411: romdata_int <= 'h412; // Line Descriptor
    6412: romdata_int <= 'h0;
    6413: romdata_int <= 'h6b0;
    6414: romdata_int <= 'h1504;
    6415: romdata_int <= 'h412; // Line Descriptor
    6416: romdata_int <= 'h200;
    6417: romdata_int <= 'h521;
    6418: romdata_int <= 'h1075;
    6419: romdata_int <= 'h412; // Line Descriptor
    6420: romdata_int <= 'h400;
    6421: romdata_int <= 'h1962;
    6422: romdata_int <= 'h735;
    6423: romdata_int <= 'h412; // Line Descriptor
    6424: romdata_int <= 'h600;
    6425: romdata_int <= 'h213d;
    6426: romdata_int <= 'h1661;
    6427: romdata_int <= 'h412; // Line Descriptor
    6428: romdata_int <= 'h800;
    6429: romdata_int <= 'h1e9b;
    6430: romdata_int <= 'h15c;
    6431: romdata_int <= 'h412; // Line Descriptor
    6432: romdata_int <= 'ha00;
    6433: romdata_int <= 'h1c42;
    6434: romdata_int <= 'hc91;
    6435: romdata_int <= 'h412; // Line Descriptor
    6436: romdata_int <= 'hc00;
    6437: romdata_int <= 'h1438;
    6438: romdata_int <= 'h8b4;
    6439: romdata_int <= 'h412; // Line Descriptor
    6440: romdata_int <= 'he00;
    6441: romdata_int <= 'h8df;
    6442: romdata_int <= 'h1f25;
    6443: romdata_int <= 'h412; // Line Descriptor
    6444: romdata_int <= 'h1000;
    6445: romdata_int <= 'he7d;
    6446: romdata_int <= 'heaa;
    6447: romdata_int <= 'h412; // Line Descriptor
    6448: romdata_int <= 'h1200;
    6449: romdata_int <= 'h2289;
    6450: romdata_int <= 'h1aaa;
    6451: romdata_int <= 'h412; // Line Descriptor
    6452: romdata_int <= 'h1400;
    6453: romdata_int <= 'h1042;
    6454: romdata_int <= 'h328;
    6455: romdata_int <= 'h412; // Line Descriptor
    6456: romdata_int <= 'h1600;
    6457: romdata_int <= 'h224;
    6458: romdata_int <= 'h18d9;
    6459: romdata_int <= 'h412; // Line Descriptor
    6460: romdata_int <= 'h1800;
    6461: romdata_int <= 'h16d2;
    6462: romdata_int <= 'h12fe;
    6463: romdata_int <= 'h412; // Line Descriptor
    6464: romdata_int <= 'h1a00;
    6465: romdata_int <= 'hd17;
    6466: romdata_int <= 'had3;
    6467: romdata_int <= 'h412; // Line Descriptor
    6468: romdata_int <= 'h1c00;
    6469: romdata_int <= 'haad;
    6470: romdata_int <= 'h1cc2;
    6471: romdata_int <= 'h412; // Line Descriptor
    6472: romdata_int <= 'h1e00;
    6473: romdata_int <= 'h1309;
    6474: romdata_int <= 'h2217;
    6475: romdata_int <= 'h412; // Line Descriptor
    6476: romdata_int <= 'h2000;
    6477: romdata_int <= 'hd8;
    6478: romdata_int <= 'h532;
    6479: romdata_int <= 'h412; // Line Descriptor
    6480: romdata_int <= 'h2200;
    6481: romdata_int <= 'h1af3;
    6482: romdata_int <= 'h20e2;
    6483: romdata_int <= 'h412; // Line Descriptor
    6484: romdata_int <= 'h0;
    6485: romdata_int <= 'h944;
    6486: romdata_int <= 'h5e;
    6487: romdata_int <= 'h412; // Line Descriptor
    6488: romdata_int <= 'h200;
    6489: romdata_int <= 'h1d1c;
    6490: romdata_int <= 'h203b;
    6491: romdata_int <= 'h412; // Line Descriptor
    6492: romdata_int <= 'h400;
    6493: romdata_int <= 'h1f3d;
    6494: romdata_int <= 'h1356;
    6495: romdata_int <= 'h412; // Line Descriptor
    6496: romdata_int <= 'h600;
    6497: romdata_int <= 'h18c4;
    6498: romdata_int <= 'h1e8a;
    6499: romdata_int <= 'h412; // Line Descriptor
    6500: romdata_int <= 'h800;
    6501: romdata_int <= 'h167b;
    6502: romdata_int <= 'h1960;
    6503: romdata_int <= 'h412; // Line Descriptor
    6504: romdata_int <= 'ha00;
    6505: romdata_int <= 'h3a;
    6506: romdata_int <= 'h1052;
    6507: romdata_int <= 'h412; // Line Descriptor
    6508: romdata_int <= 'hc00;
    6509: romdata_int <= 'hb5f;
    6510: romdata_int <= 'h14e0;
    6511: romdata_int <= 'h412; // Line Descriptor
    6512: romdata_int <= 'he00;
    6513: romdata_int <= 'h2248;
    6514: romdata_int <= 'hb37;
    6515: romdata_int <= 'h412; // Line Descriptor
    6516: romdata_int <= 'h1000;
    6517: romdata_int <= 'he48;
    6518: romdata_int <= 'h8c2;
    6519: romdata_int <= 'h412; // Line Descriptor
    6520: romdata_int <= 'h1200;
    6521: romdata_int <= 'hcc3;
    6522: romdata_int <= 'h6ca;
    6523: romdata_int <= 'h412; // Line Descriptor
    6524: romdata_int <= 'h1400;
    6525: romdata_int <= 'h1b1e;
    6526: romdata_int <= 'he7f;
    6527: romdata_int <= 'h412; // Line Descriptor
    6528: romdata_int <= 'h1600;
    6529: romdata_int <= 'h504;
    6530: romdata_int <= 'h16d5;
    6531: romdata_int <= 'h412; // Line Descriptor
    6532: romdata_int <= 'h1800;
    6533: romdata_int <= 'h6a9;
    6534: romdata_int <= 'h1a23;
    6535: romdata_int <= 'h412; // Line Descriptor
    6536: romdata_int <= 'h1a00;
    6537: romdata_int <= 'h149c;
    6538: romdata_int <= 'hc91;
    6539: romdata_int <= 'h412; // Line Descriptor
    6540: romdata_int <= 'h1c00;
    6541: romdata_int <= 'h12b5;
    6542: romdata_int <= 'h224;
    6543: romdata_int <= 'h412; // Line Descriptor
    6544: romdata_int <= 'h1e00;
    6545: romdata_int <= 'h115a;
    6546: romdata_int <= 'h2220;
    6547: romdata_int <= 'h412; // Line Descriptor
    6548: romdata_int <= 'h2000;
    6549: romdata_int <= 'h2023;
    6550: romdata_int <= 'h1ca3;
    6551: romdata_int <= 'h412; // Line Descriptor
    6552: romdata_int <= 'h2200;
    6553: romdata_int <= 'h2ea;
    6554: romdata_int <= 'h450;
    6555: romdata_int <= 'h412; // Line Descriptor
    6556: romdata_int <= 'h0;
    6557: romdata_int <= 'h341;
    6558: romdata_int <= 'h1858;
    6559: romdata_int <= 'h412; // Line Descriptor
    6560: romdata_int <= 'h200;
    6561: romdata_int <= 'h1285;
    6562: romdata_int <= 'h1a44;
    6563: romdata_int <= 'h412; // Line Descriptor
    6564: romdata_int <= 'h400;
    6565: romdata_int <= 'h67b;
    6566: romdata_int <= 'h454;
    6567: romdata_int <= 'h412; // Line Descriptor
    6568: romdata_int <= 'h600;
    6569: romdata_int <= 'h1737;
    6570: romdata_int <= 'h1c27;
    6571: romdata_int <= 'h412; // Line Descriptor
    6572: romdata_int <= 'h800;
    6573: romdata_int <= 'hf1e;
    6574: romdata_int <= 'hcd6;
    6575: romdata_int <= 'h412; // Line Descriptor
    6576: romdata_int <= 'ha00;
    6577: romdata_int <= 'ha54;
    6578: romdata_int <= 'h2048;
    6579: romdata_int <= 'h412; // Line Descriptor
    6580: romdata_int <= 'hc00;
    6581: romdata_int <= 'h208d;
    6582: romdata_int <= 'h10af;
    6583: romdata_int <= 'h412; // Line Descriptor
    6584: romdata_int <= 'he00;
    6585: romdata_int <= 'hd25;
    6586: romdata_int <= 'h1e92;
    6587: romdata_int <= 'h412; // Line Descriptor
    6588: romdata_int <= 'h1000;
    6589: romdata_int <= 'h915;
    6590: romdata_int <= 'h64b;
    6591: romdata_int <= 'h412; // Line Descriptor
    6592: romdata_int <= 'h1200;
    6593: romdata_int <= 'h1d39;
    6594: romdata_int <= 'h41;
    6595: romdata_int <= 'h412; // Line Descriptor
    6596: romdata_int <= 'h1400;
    6597: romdata_int <= 'h40;
    6598: romdata_int <= 'h14f2;
    6599: romdata_int <= 'h412; // Line Descriptor
    6600: romdata_int <= 'h1600;
    6601: romdata_int <= 'h1ec5;
    6602: romdata_int <= 'h92a;
    6603: romdata_int <= 'h412; // Line Descriptor
    6604: romdata_int <= 'h1800;
    6605: romdata_int <= 'h22c6;
    6606: romdata_int <= 'he4e;
    6607: romdata_int <= 'h412; // Line Descriptor
    6608: romdata_int <= 'h1a00;
    6609: romdata_int <= 'h1b39;
    6610: romdata_int <= 'h2302;
    6611: romdata_int <= 'h412; // Line Descriptor
    6612: romdata_int <= 'h1c00;
    6613: romdata_int <= 'h1855;
    6614: romdata_int <= 'h32c;
    6615: romdata_int <= 'h412; // Line Descriptor
    6616: romdata_int <= 'h1e00;
    6617: romdata_int <= 'h51a;
    6618: romdata_int <= 'ha95;
    6619: romdata_int <= 'h412; // Line Descriptor
    6620: romdata_int <= 'h2000;
    6621: romdata_int <= 'h1411;
    6622: romdata_int <= 'h1261;
    6623: romdata_int <= 'h512; // Line Descriptor
    6624: romdata_int <= 'h2200;
    6625: romdata_int <= 'h10bc;
    6626: romdata_int <= 'h166e;
    6627: romdata_int <= 'h1624; // Line Descriptor
    6628: romdata_int <= 'h3eae;
    6629: romdata_int <= 'h1d0b;
    6630: romdata_int <= 'h2008;
    6631: romdata_int <= 'h36d5;
    6632: romdata_int <= 'h1e86;
    6633: romdata_int <= 'h889;
    6634: romdata_int <= 'h82e;
    6635: romdata_int <= 'h4;
    6636: romdata_int <= 'hf37;
    6637: romdata_int <= 'h2e9a;
    6638: romdata_int <= 'h16b0;
    6639: romdata_int <= 'h3b5c;
    6640: romdata_int <= 'h1624; // Line Descriptor
    6641: romdata_int <= 'h4728;
    6642: romdata_int <= 'h288a;
    6643: romdata_int <= 'he6b;
    6644: romdata_int <= 'h3467;
    6645: romdata_int <= 'h1655;
    6646: romdata_int <= 'h461;
    6647: romdata_int <= 'h26d5;
    6648: romdata_int <= 'h231e;
    6649: romdata_int <= 'h30a5;
    6650: romdata_int <= 'hae0;
    6651: romdata_int <= 'h20e6;
    6652: romdata_int <= 'h534;
    6653: romdata_int <= 'h1624; // Line Descriptor
    6654: romdata_int <= 'h152b;
    6655: romdata_int <= 'h1a64;
    6656: romdata_int <= 'h3090;
    6657: romdata_int <= 'h2336;
    6658: romdata_int <= 'h10d5;
    6659: romdata_int <= 'h2a62;
    6660: romdata_int <= 'h44f2;
    6661: romdata_int <= 'h3eb6;
    6662: romdata_int <= 'h6c9;
    6663: romdata_int <= 'h3354;
    6664: romdata_int <= 'h144a;
    6665: romdata_int <= 'h1077;
    6666: romdata_int <= 'h1624; // Line Descriptor
    6667: romdata_int <= 'h3349;
    6668: romdata_int <= 'h67;
    6669: romdata_int <= 'haa6;
    6670: romdata_int <= 'hcf2;
    6671: romdata_int <= 'h1888;
    6672: romdata_int <= 'h3d27;
    6673: romdata_int <= 'h2bd;
    6674: romdata_int <= 'h2c5c;
    6675: romdata_int <= 'h4648;
    6676: romdata_int <= 'h2b22;
    6677: romdata_int <= 'h4301;
    6678: romdata_int <= 'h4134;
    6679: romdata_int <= 'h424; // Line Descriptor
    6680: romdata_int <= 'h40d9;
    6681: romdata_int <= 'h2655;
    6682: romdata_int <= 'h132b;
    6683: romdata_int <= 'h424; // Line Descriptor
    6684: romdata_int <= 'h25e;
    6685: romdata_int <= 'h252d;
    6686: romdata_int <= 'h2e9f;
    6687: romdata_int <= 'h424; // Line Descriptor
    6688: romdata_int <= 'h3825;
    6689: romdata_int <= 'h2d4d;
    6690: romdata_int <= 'h4552;
    6691: romdata_int <= 'h424; // Line Descriptor
    6692: romdata_int <= 'h42ab;
    6693: romdata_int <= 'h3a75;
    6694: romdata_int <= 'h641;
    6695: romdata_int <= 'h524; // Line Descriptor
    6696: romdata_int <= 'h1911;
    6697: romdata_int <= 'h2561;
    6698: romdata_int <= 'h128a;
    6699: romdata_int <= 'h161e; // Line Descriptor
    6700: romdata_int <= 'h340d;
    6701: romdata_int <= 'h3b28;
    6702: romdata_int <= 'h208a;
    6703: romdata_int <= 'hc6b;
    6704: romdata_int <= 'h2c67;
    6705: romdata_int <= 'h1455;
    6706: romdata_int <= 'h461;
    6707: romdata_int <= 'h1ed5;
    6708: romdata_int <= 'h1b1e;
    6709: romdata_int <= 'h26a5;
    6710: romdata_int <= 'h6e0;
    6711: romdata_int <= 'h18e6;
    6712: romdata_int <= 'h161e; // Line Descriptor
    6713: romdata_int <= 'h112b;
    6714: romdata_int <= 'h1664;
    6715: romdata_int <= 'h2690;
    6716: romdata_int <= 'h1936;
    6717: romdata_int <= 'hcd5;
    6718: romdata_int <= 'h2262;
    6719: romdata_int <= 'h38f2;
    6720: romdata_int <= 'h32b6;
    6721: romdata_int <= 'h2c9;
    6722: romdata_int <= 'h2554;
    6723: romdata_int <= 'hc4a;
    6724: romdata_int <= 'ha77;
    6725: romdata_int <= 'h161e; // Line Descriptor
    6726: romdata_int <= 'h2e70;
    6727: romdata_int <= 'h134f;
    6728: romdata_int <= 'h825;
    6729: romdata_int <= 'h254d;
    6730: romdata_int <= 'hf52;
    6731: romdata_int <= 'h3138;
    6732: romdata_int <= 'h8f;
    6733: romdata_int <= 'h1c0e;
    6734: romdata_int <= 'h12ab;
    6735: romdata_int <= 'h3475;
    6736: romdata_int <= 'h1e41;
    6737: romdata_int <= 'h164c;
    6738: romdata_int <= 'h161e; // Line Descriptor
    6739: romdata_int <= 'he5d;
    6740: romdata_int <= 'h67b;
    6741: romdata_int <= 'h32fd;
    6742: romdata_int <= 'h36eb;
    6743: romdata_int <= 'h2e18;
    6744: romdata_int <= 'h2a40;
    6745: romdata_int <= 'h2122;
    6746: romdata_int <= 'hacf;
    6747: romdata_int <= 'h80;
    6748: romdata_int <= 'h14ab;
    6749: romdata_int <= 'h2c98;
    6750: romdata_int <= 'h28b4;
    6751: romdata_int <= 'h161e; // Line Descriptor
    6752: romdata_int <= 'h28cb;
    6753: romdata_int <= 'h31d;
    6754: romdata_int <= 'h1e32;
    6755: romdata_int <= 'h30f6;
    6756: romdata_int <= 'h26a2;
    6757: romdata_int <= 'h34a4;
    6758: romdata_int <= 'h1ab3;
    6759: romdata_int <= 'h23d;
    6760: romdata_int <= 'h2a72;
    6761: romdata_int <= 'h3b3e;
    6762: romdata_int <= 'h55d;
    6763: romdata_int <= 'h208f;
    6764: romdata_int <= 'h41e; // Line Descriptor
    6765: romdata_int <= 'ha32;
    6766: romdata_int <= 'h18bd;
    6767: romdata_int <= 'h1103;
    6768: romdata_int <= 'h41e; // Line Descriptor
    6769: romdata_int <= 'h4ef;
    6770: romdata_int <= 'h28e3;
    6771: romdata_int <= 'h2edc;
    6772: romdata_int <= 'h41e; // Line Descriptor
    6773: romdata_int <= 'h2af2;
    6774: romdata_int <= 'h1683;
    6775: romdata_int <= 'h3274;
    6776: romdata_int <= 'h41e; // Line Descriptor
    6777: romdata_int <= 'h1556;
    6778: romdata_int <= 'h3b20;
    6779: romdata_int <= 'h1c1e;
    6780: romdata_int <= 'h41e; // Line Descriptor
    6781: romdata_int <= 'h2c78;
    6782: romdata_int <= 'h6fc;
    6783: romdata_int <= 'h3938;
    6784: romdata_int <= 'h41e; // Line Descriptor
    6785: romdata_int <= 'h14b;
    6786: romdata_int <= 'h24a8;
    6787: romdata_int <= 'h3097;
    6788: romdata_int <= 'h41e; // Line Descriptor
    6789: romdata_int <= 'h1ca1;
    6790: romdata_int <= 'h1340;
    6791: romdata_int <= 'he5a;
    6792: romdata_int <= 'h41e; // Line Descriptor
    6793: romdata_int <= 'h1ae5;
    6794: romdata_int <= 'h366b;
    6795: romdata_int <= 'h839;
    6796: romdata_int <= 'h41e; // Line Descriptor
    6797: romdata_int <= 'h389e;
    6798: romdata_int <= 'h1081;
    6799: romdata_int <= 'h374d;
    6800: romdata_int <= 'h51e; // Line Descriptor
    6801: romdata_int <= 'h2351;
    6802: romdata_int <= 'h86f;
    6803: romdata_int <= 'h2313;
    6804: romdata_int <= 'h161b; // Line Descriptor
    6805: romdata_int <= 'hed1;
    6806: romdata_int <= 'h1899;
    6807: romdata_int <= 'h544;
    6808: romdata_int <= 'h2015;
    6809: romdata_int <= 'h30f8;
    6810: romdata_int <= 'h332a;
    6811: romdata_int <= 'h1c17;
    6812: romdata_int <= 'h1841;
    6813: romdata_int <= 'h2a31;
    6814: romdata_int <= 'h1500;
    6815: romdata_int <= 'h121b;
    6816: romdata_int <= 'h20f6;
    6817: romdata_int <= 'h161b; // Line Descriptor
    6818: romdata_int <= 'h34d2;
    6819: romdata_int <= 'h163e;
    6820: romdata_int <= 'h2a76;
    6821: romdata_int <= 'h140f;
    6822: romdata_int <= 'h3503;
    6823: romdata_int <= 'h2ba;
    6824: romdata_int <= 'h26cf;
    6825: romdata_int <= 'h1a60;
    6826: romdata_int <= 'h281f;
    6827: romdata_int <= 'h700;
    6828: romdata_int <= 'h1e41;
    6829: romdata_int <= 'h3128;
    6830: romdata_int <= 'h161b; // Line Descriptor
    6831: romdata_int <= 'h2e93;
    6832: romdata_int <= 'h1e1c;
    6833: romdata_int <= 'h651;
    6834: romdata_int <= 'h2d0c;
    6835: romdata_int <= 'hd4c;
    6836: romdata_int <= 'h2120;
    6837: romdata_int <= 'h2842;
    6838: romdata_int <= 'h645;
    6839: romdata_int <= 'h10e3;
    6840: romdata_int <= 'h1947;
    6841: romdata_int <= 'h2c20;
    6842: romdata_int <= 'h1c47;
    6843: romdata_int <= 'h161b; // Line Descriptor
    6844: romdata_int <= 'h898;
    6845: romdata_int <= 'h28c;
    6846: romdata_int <= 'h2318;
    6847: romdata_int <= 'hcfc;
    6848: romdata_int <= 'hf59;
    6849: romdata_int <= 'h2530;
    6850: romdata_int <= 'h2ec7;
    6851: romdata_int <= 'h10d9;
    6852: romdata_int <= 'ha4;
    6853: romdata_int <= 'h3346;
    6854: romdata_int <= 'h231f;
    6855: romdata_int <= 'h1a53;
    6856: romdata_int <= 'h161b; // Line Descriptor
    6857: romdata_int <= 'h109d;
    6858: romdata_int <= 'h3020;
    6859: romdata_int <= 'h28a1;
    6860: romdata_int <= 'h2746;
    6861: romdata_int <= 'h2b65;
    6862: romdata_int <= 'hc;
    6863: romdata_int <= 'had9;
    6864: romdata_int <= 'h2cb0;
    6865: romdata_int <= 'h1608;
    6866: romdata_int <= 'hb24;
    6867: romdata_int <= 'hced;
    6868: romdata_int <= 'h354b;
    6869: romdata_int <= 'h161b; // Line Descriptor
    6870: romdata_int <= 'h167;
    6871: romdata_int <= 'h1c12;
    6872: romdata_int <= 'h125d;
    6873: romdata_int <= 'h1a52;
    6874: romdata_int <= 'h443;
    6875: romdata_int <= 'h1f59;
    6876: romdata_int <= 'h1647;
    6877: romdata_int <= 'h14be;
    6878: romdata_int <= 'he95;
    6879: romdata_int <= 'h24b2;
    6880: romdata_int <= 'h2e1d;
    6881: romdata_int <= 'h474;
    6882: romdata_int <= 'h41b; // Line Descriptor
    6883: romdata_int <= 'ha3d;
    6884: romdata_int <= 'h232e;
    6885: romdata_int <= 'h835;
    6886: romdata_int <= 'h41b; // Line Descriptor
    6887: romdata_int <= 'h247c;
    6888: romdata_int <= 'h12f2;
    6889: romdata_int <= 'h268a;
    6890: romdata_int <= 'h41b; // Line Descriptor
    6891: romdata_int <= 'h3357;
    6892: romdata_int <= 'h93b;
    6893: romdata_int <= 'h2ac;
    6894: romdata_int <= 'h41b; // Line Descriptor
    6895: romdata_int <= 'h3511;
    6896: romdata_int <= 'h18d6;
    6897: romdata_int <= 'h114c;
    6898: romdata_int <= 'h41b; // Line Descriptor
    6899: romdata_int <= 'h12f4;
    6900: romdata_int <= 'h2aa3;
    6901: romdata_int <= 'h2242;
    6902: romdata_int <= 'h41b; // Line Descriptor
    6903: romdata_int <= 'h1f57;
    6904: romdata_int <= 'h2495;
    6905: romdata_int <= 'h1a8e;
    6906: romdata_int <= 'h41b; // Line Descriptor
    6907: romdata_int <= 'h2141;
    6908: romdata_int <= 'hf11;
    6909: romdata_int <= 'hab7;
    6910: romdata_int <= 'h41b; // Line Descriptor
    6911: romdata_int <= 'h4c6;
    6912: romdata_int <= 'h2c49;
    6913: romdata_int <= 'hd54;
    6914: romdata_int <= 'h41b; // Line Descriptor
    6915: romdata_int <= 'h2f9;
    6916: romdata_int <= 'h314d;
    6917: romdata_int <= 'h6d1;
    6918: romdata_int <= 'h41b; // Line Descriptor
    6919: romdata_int <= 'h28a6;
    6920: romdata_int <= 'h16a4;
    6921: romdata_int <= 'h2f39;
    6922: romdata_int <= 'h41b; // Line Descriptor
    6923: romdata_int <= 'h8bd;
    6924: romdata_int <= 'h330f;
    6925: romdata_int <= 'h275d;
    6926: romdata_int <= 'h51b; // Line Descriptor
    6927: romdata_int <= 'h1433;
    6928: romdata_int <= 'h14a;
    6929: romdata_int <= 'h1c62;
    6930: romdata_int <= 'he19; // Line Descriptor
    6931: romdata_int <= 'h2800;
    6932: romdata_int <= 'h181c;
    6933: romdata_int <= 'h165f;
    6934: romdata_int <= 'h8fe;
    6935: romdata_int <= 'h16a2;
    6936: romdata_int <= 'h182a;
    6937: romdata_int <= 'h28c9;
    6938: romdata_int <= 'h10ce;
    6939: romdata_int <= 'he19; // Line Descriptor
    6940: romdata_int <= 'h2a00;
    6941: romdata_int <= 'h2465;
    6942: romdata_int <= 'h2ee5;
    6943: romdata_int <= 'h2cc0;
    6944: romdata_int <= 'h2e5d;
    6945: romdata_int <= 'h1c7b;
    6946: romdata_int <= 'h6fd;
    6947: romdata_int <= 'h2eb;
    6948: romdata_int <= 'he19; // Line Descriptor
    6949: romdata_int <= 'h2c00;
    6950: romdata_int <= 'h225;
    6951: romdata_int <= 'h2e4;
    6952: romdata_int <= 'h260a;
    6953: romdata_int <= 'h2493;
    6954: romdata_int <= 'h1a61;
    6955: romdata_int <= 'h1e7f;
    6956: romdata_int <= 'he8c;
    6957: romdata_int <= 'he19; // Line Descriptor
    6958: romdata_int <= 'h2e00;
    6959: romdata_int <= 'h470;
    6960: romdata_int <= 'h28b4;
    6961: romdata_int <= 'h48f;
    6962: romdata_int <= 'h30d4;
    6963: romdata_int <= 'h202b;
    6964: romdata_int <= 'h22ba;
    6965: romdata_int <= 'h30b1;
    6966: romdata_int <= 'he19; // Line Descriptor
    6967: romdata_int <= 'h3000;
    6968: romdata_int <= 'h1ecd;
    6969: romdata_int <= 'h650;
    6970: romdata_int <= 'h1a32;
    6971: romdata_int <= 'h22bd;
    6972: romdata_int <= 'h2d03;
    6973: romdata_int <= 'h142f;
    6974: romdata_int <= 'h4f8;
    6975: romdata_int <= 'h419; // Line Descriptor
    6976: romdata_int <= 'h0;
    6977: romdata_int <= 'h2aa1;
    6978: romdata_int <= 'h1315;
    6979: romdata_int <= 'h419; // Line Descriptor
    6980: romdata_int <= 'h200;
    6981: romdata_int <= 'ha72;
    6982: romdata_int <= 'h2002;
    6983: romdata_int <= 'h419; // Line Descriptor
    6984: romdata_int <= 'h400;
    6985: romdata_int <= 'h270b;
    6986: romdata_int <= 'h1808;
    6987: romdata_int <= 'h419; // Line Descriptor
    6988: romdata_int <= 'h600;
    6989: romdata_int <= 'h1c89;
    6990: romdata_int <= 'h102e;
    6991: romdata_int <= 'h419; // Line Descriptor
    6992: romdata_int <= 'h800;
    6993: romdata_int <= 'h9a;
    6994: romdata_int <= 'h2cb0;
    6995: romdata_int <= 'h419; // Line Descriptor
    6996: romdata_int <= 'ha00;
    6997: romdata_int <= 'h30ec;
    6998: romdata_int <= 'h1e0b;
    6999: romdata_int <= 'h419; // Line Descriptor
    7000: romdata_int <= 'hc00;
    7001: romdata_int <= 'h223a;
    7002: romdata_int <= 'h30a1;
    7003: romdata_int <= 'h419; // Line Descriptor
    7004: romdata_int <= 'he00;
    7005: romdata_int <= 'h2938;
    7006: romdata_int <= 'h2259;
    7007: romdata_int <= 'h419; // Line Descriptor
    7008: romdata_int <= 'h1000;
    7009: romdata_int <= 'hcb8;
    7010: romdata_int <= 'ha7b;
    7011: romdata_int <= 'h419; // Line Descriptor
    7012: romdata_int <= 'h1200;
    7013: romdata_int <= 'h10b9;
    7014: romdata_int <= 'h53b;
    7015: romdata_int <= 'h419; // Line Descriptor
    7016: romdata_int <= 'h1400;
    7017: romdata_int <= 'h129b;
    7018: romdata_int <= 'h2512;
    7019: romdata_int <= 'h419; // Line Descriptor
    7020: romdata_int <= 'h1600;
    7021: romdata_int <= 'h1565;
    7022: romdata_int <= 'h2ac7;
    7023: romdata_int <= 'h419; // Line Descriptor
    7024: romdata_int <= 'h1800;
    7025: romdata_int <= 'h679;
    7026: romdata_int <= 'h1c1e;
    7027: romdata_int <= 'h419; // Line Descriptor
    7028: romdata_int <= 'h1a00;
    7029: romdata_int <= 'h1aef;
    7030: romdata_int <= 'he2a;
    7031: romdata_int <= 'h519; // Line Descriptor
    7032: romdata_int <= 'h1c00;
    7033: romdata_int <= 'h1728;
    7034: romdata_int <= 'h8a;
    7035: romdata_int <= 'h1612; // Line Descriptor
    7036: romdata_int <= 'h1699;
    7037: romdata_int <= 'hf3d;
    7038: romdata_int <= 'h165;
    7039: romdata_int <= 'h1cc7;
    7040: romdata_int <= 'hc4c;
    7041: romdata_int <= 'hb0b;
    7042: romdata_int <= 'h879;
    7043: romdata_int <= 'h81e;
    7044: romdata_int <= 'h14bc;
    7045: romdata_int <= 'h1c9d;
    7046: romdata_int <= 'h10ef;
    7047: romdata_int <= 'h1e2a;
    7048: romdata_int <= 'h1612; // Line Descriptor
    7049: romdata_int <= 'h313;
    7050: romdata_int <= 'h1a0b;
    7051: romdata_int <= 'h187a;
    7052: romdata_int <= 'h628;
    7053: romdata_int <= 'h845;
    7054: romdata_int <= 'h18a2;
    7055: romdata_int <= 'h416;
    7056: romdata_int <= 'h1f3e;
    7057: romdata_int <= 'h1a0e;
    7058: romdata_int <= 'h737;
    7059: romdata_int <= 'h234c;
    7060: romdata_int <= 'ha91;
    7061: romdata_int <= 'h1612; // Line Descriptor
    7062: romdata_int <= 'h180b;
    7063: romdata_int <= 'h1d06;
    7064: romdata_int <= 'h2340;
    7065: romdata_int <= 'hac;
    7066: romdata_int <= 'h20ed;
    7067: romdata_int <= 'h155a;
    7068: romdata_int <= 'hf12;
    7069: romdata_int <= 'h63e;
    7070: romdata_int <= 'h367;
    7071: romdata_int <= 'hd26;
    7072: romdata_int <= 'h55f;
    7073: romdata_int <= 'h4df;
    7074: romdata_int <= 'h1612; // Line Descriptor
    7075: romdata_int <= 'h12e7;
    7076: romdata_int <= 'h1672;
    7077: romdata_int <= 'hb08;
    7078: romdata_int <= 'heaf;
    7079: romdata_int <= 'h193a;
    7080: romdata_int <= 'h1cdb;
    7081: romdata_int <= 'h1f4f;
    7082: romdata_int <= 'ha1f;
    7083: romdata_int <= 'hee;
    7084: romdata_int <= 'h1687;
    7085: romdata_int <= 'h14bd;
    7086: romdata_int <= 'h215f;
    7087: romdata_int <= 'h1612; // Line Descriptor
    7088: romdata_int <= 'hee9;
    7089: romdata_int <= 'h2086;
    7090: romdata_int <= 'h14f8;
    7091: romdata_int <= 'ha03;
    7092: romdata_int <= 'h165f;
    7093: romdata_int <= 'h2028;
    7094: romdata_int <= 'h12a6;
    7095: romdata_int <= 'h1c17;
    7096: romdata_int <= 'h12d3;
    7097: romdata_int <= 'h254;
    7098: romdata_int <= 'h2106;
    7099: romdata_int <= 'h758;
    7100: romdata_int <= 'h1612; // Line Descriptor
    7101: romdata_int <= 'hc94;
    7102: romdata_int <= 'h6ab;
    7103: romdata_int <= 'h131d;
    7104: romdata_int <= 'h14cf;
    7105: romdata_int <= 'h26f;
    7106: romdata_int <= 'h747;
    7107: romdata_int <= 'hcf2;
    7108: romdata_int <= 'h10d3;
    7109: romdata_int <= 'h20fb;
    7110: romdata_int <= 'h132c;
    7111: romdata_int <= 'h1962;
    7112: romdata_int <= 'h1b42;
    7113: romdata_int <= 'h1612; // Line Descriptor
    7114: romdata_int <= 'h1132;
    7115: romdata_int <= 'h45a;
    7116: romdata_int <= 'h10a1;
    7117: romdata_int <= 'h12b6;
    7118: romdata_int <= 'h1e45;
    7119: romdata_int <= 'h342;
    7120: romdata_int <= 'hd4;
    7121: romdata_int <= 'he2d;
    7122: romdata_int <= 'h1630;
    7123: romdata_int <= 'he80;
    7124: romdata_int <= 'h1ec4;
    7125: romdata_int <= 'h2242;
    7126: romdata_int <= 'h1612; // Line Descriptor
    7127: romdata_int <= 'h1ceb;
    7128: romdata_int <= 'hc79;
    7129: romdata_int <= 'h1f2c;
    7130: romdata_int <= 'h1a5e;
    7131: romdata_int <= 'h1139;
    7132: romdata_int <= 'h110f;
    7133: romdata_int <= 'h1681;
    7134: romdata_int <= 'h220f;
    7135: romdata_int <= 'h1866;
    7136: romdata_int <= 'ha3e;
    7137: romdata_int <= 'h1ac7;
    7138: romdata_int <= 'h154e;
    7139: romdata_int <= 'h1612; // Line Descriptor
    7140: romdata_int <= 'h77;
    7141: romdata_int <= 'h89d;
    7142: romdata_int <= 'h2e2;
    7143: romdata_int <= 'h53a;
    7144: romdata_int <= 'h2247;
    7145: romdata_int <= 'h22a3;
    7146: romdata_int <= 'h1ad9;
    7147: romdata_int <= 'hc4b;
    7148: romdata_int <= 'h431;
    7149: romdata_int <= 'h863;
    7150: romdata_int <= 'h16;
    7151: romdata_int <= 'h907;
    7152: romdata_int <= 'h412; // Line Descriptor
    7153: romdata_int <= 'h0;
    7154: romdata_int <= 'h278;
    7155: romdata_int <= 'he93;
    7156: romdata_int <= 'h412; // Line Descriptor
    7157: romdata_int <= 'h200;
    7158: romdata_int <= 'h184c;
    7159: romdata_int <= 'h651;
    7160: romdata_int <= 'h412; // Line Descriptor
    7161: romdata_int <= 'h400;
    7162: romdata_int <= 'h8b;
    7163: romdata_int <= 'h22cd;
    7164: romdata_int <= 'h412; // Line Descriptor
    7165: romdata_int <= 'h600;
    7166: romdata_int <= 'h16dc;
    7167: romdata_int <= 'h1a3a;
    7168: romdata_int <= 'h412; // Line Descriptor
    7169: romdata_int <= 'h800;
    7170: romdata_int <= 'h134c;
    7171: romdata_int <= 'h1d50;
    7172: romdata_int <= 'h412; // Line Descriptor
    7173: romdata_int <= 'ha00;
    7174: romdata_int <= 'ha60;
    7175: romdata_int <= 'h214e;
    7176: romdata_int <= 'h412; // Line Descriptor
    7177: romdata_int <= 'hc00;
    7178: romdata_int <= 'hcd2;
    7179: romdata_int <= 'h146b;
    7180: romdata_int <= 'h412; // Line Descriptor
    7181: romdata_int <= 'he00;
    7182: romdata_int <= 'h10ee;
    7183: romdata_int <= 'h435;
    7184: romdata_int <= 'h412; // Line Descriptor
    7185: romdata_int <= 'h1000;
    7186: romdata_int <= 'h93c;
    7187: romdata_int <= 'h1ebd;
    7188: romdata_int <= 'h412; // Line Descriptor
    7189: romdata_int <= 'h1200;
    7190: romdata_int <= 'h1c0e;
    7191: romdata_int <= 'h10f;
    7192: romdata_int <= 'h412; // Line Descriptor
    7193: romdata_int <= 'h1400;
    7194: romdata_int <= 'h2310;
    7195: romdata_int <= 'heb4;
    7196: romdata_int <= 'h412; // Line Descriptor
    7197: romdata_int <= 'h1600;
    7198: romdata_int <= 'h1708;
    7199: romdata_int <= 'h1ada;
    7200: romdata_int <= 'h412; // Line Descriptor
    7201: romdata_int <= 'h1800;
    7202: romdata_int <= 'h10c7;
    7203: romdata_int <= 'haa1;
    7204: romdata_int <= 'h412; // Line Descriptor
    7205: romdata_int <= 'h1a00;
    7206: romdata_int <= 'h148e;
    7207: romdata_int <= 'h6ea;
    7208: romdata_int <= 'h412; // Line Descriptor
    7209: romdata_int <= 'h1c00;
    7210: romdata_int <= 'hd21;
    7211: romdata_int <= 'h1305;
    7212: romdata_int <= 'h412; // Line Descriptor
    7213: romdata_int <= 'h1e00;
    7214: romdata_int <= 'h20da;
    7215: romdata_int <= 'h8bc;
    7216: romdata_int <= 'h412; // Line Descriptor
    7217: romdata_int <= 'h2000;
    7218: romdata_int <= 'h1f1b;
    7219: romdata_int <= 'h4fd;
    7220: romdata_int <= 'h512; // Line Descriptor
    7221: romdata_int <= 'h2200;
    7222: romdata_int <= 'h1910;
    7223: romdata_int <= 'h2e8;
    7224: romdata_int <= 'h180f; // Line Descriptor
    7225: romdata_int <= 'h0;
    7226: romdata_int <= 'h1c8a;
    7227: romdata_int <= 'h106b;
    7228: romdata_int <= 'h667;
    7229: romdata_int <= 'h1655;
    7230: romdata_int <= 'ha61;
    7231: romdata_int <= 'h2d5;
    7232: romdata_int <= 'hf1e;
    7233: romdata_int <= 'hca5;
    7234: romdata_int <= 'h12e0;
    7235: romdata_int <= 'h2e6;
    7236: romdata_int <= 'h134;
    7237: romdata_int <= 'h18ae;
    7238: romdata_int <= 'h180f; // Line Descriptor
    7239: romdata_int <= 'h200;
    7240: romdata_int <= 'h408;
    7241: romdata_int <= 'h265;
    7242: romdata_int <= 'h1ae5;
    7243: romdata_int <= 'hc0;
    7244: romdata_int <= 'h185d;
    7245: romdata_int <= 'h47b;
    7246: romdata_int <= 'h8fd;
    7247: romdata_int <= 'h8eb;
    7248: romdata_int <= 'h1a18;
    7249: romdata_int <= 'h1640;
    7250: romdata_int <= 'h1122;
    7251: romdata_int <= 'h6cf;
    7252: romdata_int <= 'h180f; // Line Descriptor
    7253: romdata_int <= 'h400;
    7254: romdata_int <= 'h811;
    7255: romdata_int <= 'h12e2;
    7256: romdata_int <= 'h1c3d;
    7257: romdata_int <= 'h14b0;
    7258: romdata_int <= 'h1239;
    7259: romdata_int <= 'hd0a;
    7260: romdata_int <= 'h10ff;
    7261: romdata_int <= 'h407;
    7262: romdata_int <= 'hf60;
    7263: romdata_int <= 'h1c0a;
    7264: romdata_int <= 'had0;
    7265: romdata_int <= 'h149c;
    7266: romdata_int <= 'h40f; // Line Descriptor
    7267: romdata_int <= 'h600;
    7268: romdata_int <= 'h1816;
    7269: romdata_int <= 'h8eb;
    7270: romdata_int <= 'h40f; // Line Descriptor
    7271: romdata_int <= 'h800;
    7272: romdata_int <= 'h1b17;
    7273: romdata_int <= 'h48f;
    7274: romdata_int <= 'h40f; // Line Descriptor
    7275: romdata_int <= 'ha00;
    7276: romdata_int <= 'ha7d;
    7277: romdata_int <= 'hd42;
    7278: romdata_int <= 'h40f; // Line Descriptor
    7279: romdata_int <= 'hc00;
    7280: romdata_int <= 'h1301;
    7281: romdata_int <= 'hb47;
    7282: romdata_int <= 'h40f; // Line Descriptor
    7283: romdata_int <= 'he00;
    7284: romdata_int <= 'h610;
    7285: romdata_int <= 'h1866;
    7286: romdata_int <= 'h40f; // Line Descriptor
    7287: romdata_int <= 'h1000;
    7288: romdata_int <= 'h16c8;
    7289: romdata_int <= 'h165f;
    7290: romdata_int <= 'h40f; // Line Descriptor
    7291: romdata_int <= 'h1200;
    7292: romdata_int <= 'he90;
    7293: romdata_int <= 'hea7;
    7294: romdata_int <= 'h40f; // Line Descriptor
    7295: romdata_int <= 'h1400;
    7296: romdata_int <= 'h333;
    7297: romdata_int <= 'h1a42;
    7298: romdata_int <= 'h40f; // Line Descriptor
    7299: romdata_int <= 'h1600;
    7300: romdata_int <= 'hbd;
    7301: romdata_int <= 'h2f;
    7302: romdata_int <= 'h40f; // Line Descriptor
    7303: romdata_int <= 'h1800;
    7304: romdata_int <= 'hce4;
    7305: romdata_int <= 'h149d;
    7306: romdata_int <= 'h40f; // Line Descriptor
    7307: romdata_int <= 'h1a00;
    7308: romdata_int <= 'h1100;
    7309: romdata_int <= 'h1ca4;
    7310: romdata_int <= 'h40f; // Line Descriptor
    7311: romdata_int <= 'h1c00;
    7312: romdata_int <= 'h145a;
    7313: romdata_int <= 'h674;
    7314: romdata_int <= 'h40f; // Line Descriptor
    7315: romdata_int <= 'h0;
    7316: romdata_int <= 'h1a0a;
    7317: romdata_int <= 'h2a9;
    7318: romdata_int <= 'h40f; // Line Descriptor
    7319: romdata_int <= 'h200;
    7320: romdata_int <= 'h6ac;
    7321: romdata_int <= 'h144e;
    7322: romdata_int <= 'h40f; // Line Descriptor
    7323: romdata_int <= 'h400;
    7324: romdata_int <= 'h1866;
    7325: romdata_int <= 'h1c21;
    7326: romdata_int <= 'h40f; // Line Descriptor
    7327: romdata_int <= 'h600;
    7328: romdata_int <= 'h1126;
    7329: romdata_int <= 'h43;
    7330: romdata_int <= 'h40f; // Line Descriptor
    7331: romdata_int <= 'h800;
    7332: romdata_int <= 'hf5b;
    7333: romdata_int <= 'h555;
    7334: romdata_int <= 'h40f; // Line Descriptor
    7335: romdata_int <= 'ha00;
    7336: romdata_int <= 'h148f;
    7337: romdata_int <= 'h18c2;
    7338: romdata_int <= 'h40f; // Line Descriptor
    7339: romdata_int <= 'hc00;
    7340: romdata_int <= 'h417;
    7341: romdata_int <= 'h16b3;
    7342: romdata_int <= 'h40f; // Line Descriptor
    7343: romdata_int <= 'he00;
    7344: romdata_int <= 'h20f;
    7345: romdata_int <= 'hd1e;
    7346: romdata_int <= 'h40f; // Line Descriptor
    7347: romdata_int <= 'h1000;
    7348: romdata_int <= 'h68;
    7349: romdata_int <= 'he20;
    7350: romdata_int <= 'h40f; // Line Descriptor
    7351: romdata_int <= 'h1200;
    7352: romdata_int <= 'h1705;
    7353: romdata_int <= 'ha6d;
    7354: romdata_int <= 'h40f; // Line Descriptor
    7355: romdata_int <= 'h1400;
    7356: romdata_int <= 'h1c09;
    7357: romdata_int <= 'h6c3;
    7358: romdata_int <= 'h40f; // Line Descriptor
    7359: romdata_int <= 'h1600;
    7360: romdata_int <= 'h129d;
    7361: romdata_int <= 'h1025;
    7362: romdata_int <= 'h40f; // Line Descriptor
    7363: romdata_int <= 'h1800;
    7364: romdata_int <= 'ha2a;
    7365: romdata_int <= 'h1a2d;
    7366: romdata_int <= 'h40f; // Line Descriptor
    7367: romdata_int <= 'h1a00;
    7368: romdata_int <= 'hc0f;
    7369: romdata_int <= 'h870;
    7370: romdata_int <= 'h50f; // Line Descriptor
    7371: romdata_int <= 'h1c00;
    7372: romdata_int <= 'h84b;
    7373: romdata_int <= 'h1303;
    7374: romdata_int <= 'h160c; // Line Descriptor
    7375: romdata_int <= 'h600;
    7376: romdata_int <= 'hd0a;
    7377: romdata_int <= 'h1427;
    7378: romdata_int <= 'hf5e;
    7379: romdata_int <= 'ha7b;
    7380: romdata_int <= 'h254;
    7381: romdata_int <= 'hda;
    7382: romdata_int <= 'h8a0;
    7383: romdata_int <= 'hb1e;
    7384: romdata_int <= 'h42e;
    7385: romdata_int <= 'h1638;
    7386: romdata_int <= 'h296;
    7387: romdata_int <= 'h40c; // Line Descriptor
    7388: romdata_int <= 'h800;
    7389: romdata_int <= 'hadf;
    7390: romdata_int <= 'h16b1;
    7391: romdata_int <= 'h40c; // Line Descriptor
    7392: romdata_int <= 'ha00;
    7393: romdata_int <= 'h1702;
    7394: romdata_int <= 'hf4f;
    7395: romdata_int <= 'h40c; // Line Descriptor
    7396: romdata_int <= 'hc00;
    7397: romdata_int <= 'h12db;
    7398: romdata_int <= 'h319;
    7399: romdata_int <= 'h40c; // Line Descriptor
    7400: romdata_int <= 'he00;
    7401: romdata_int <= 'h53f;
    7402: romdata_int <= 'hb1f;
    7403: romdata_int <= 'h40c; // Line Descriptor
    7404: romdata_int <= 'h1000;
    7405: romdata_int <= 'h358;
    7406: romdata_int <= 'h10ab;
    7407: romdata_int <= 'h40c; // Line Descriptor
    7408: romdata_int <= 'h1200;
    7409: romdata_int <= 'h115c;
    7410: romdata_int <= 'hce4;
    7411: romdata_int <= 'h40c; // Line Descriptor
    7412: romdata_int <= 'h1400;
    7413: romdata_int <= 'h1548;
    7414: romdata_int <= 'h459;
    7415: romdata_int <= 'h40c; // Line Descriptor
    7416: romdata_int <= 'h1600;
    7417: romdata_int <= 'heba;
    7418: romdata_int <= 'h52;
    7419: romdata_int <= 'h40c; // Line Descriptor
    7420: romdata_int <= 'h0;
    7421: romdata_int <= 'hc79;
    7422: romdata_int <= 'hefc;
    7423: romdata_int <= 'h40c; // Line Descriptor
    7424: romdata_int <= 'h200;
    7425: romdata_int <= 'h6fa;
    7426: romdata_int <= 'h106e;
    7427: romdata_int <= 'h40c; // Line Descriptor
    7428: romdata_int <= 'h400;
    7429: romdata_int <= 'h125e;
    7430: romdata_int <= 'h8f;
    7431: romdata_int <= 'h40c; // Line Descriptor
    7432: romdata_int <= 'h600;
    7433: romdata_int <= 'hb;
    7434: romdata_int <= 'hb36;
    7435: romdata_int <= 'h40c; // Line Descriptor
    7436: romdata_int <= 'h800;
    7437: romdata_int <= 'ha97;
    7438: romdata_int <= 'h435;
    7439: romdata_int <= 'h40c; // Line Descriptor
    7440: romdata_int <= 'ha00;
    7441: romdata_int <= 'h1493;
    7442: romdata_int <= 'h71f;
    7443: romdata_int <= 'h40c; // Line Descriptor
    7444: romdata_int <= 'hc00;
    7445: romdata_int <= 'h112e;
    7446: romdata_int <= 'h1268;
    7447: romdata_int <= 'h40c; // Line Descriptor
    7448: romdata_int <= 'he00;
    7449: romdata_int <= 'h42d;
    7450: romdata_int <= 'h1533;
    7451: romdata_int <= 'h40c; // Line Descriptor
    7452: romdata_int <= 'h1000;
    7453: romdata_int <= 'he54;
    7454: romdata_int <= 'h2a2;
    7455: romdata_int <= 'h40c; // Line Descriptor
    7456: romdata_int <= 'h1200;
    7457: romdata_int <= 'h8a2;
    7458: romdata_int <= 'h822;
    7459: romdata_int <= 'h40c; // Line Descriptor
    7460: romdata_int <= 'h1400;
    7461: romdata_int <= 'h1652;
    7462: romdata_int <= 'hcba;
    7463: romdata_int <= 'h40c; // Line Descriptor
    7464: romdata_int <= 'h1600;
    7465: romdata_int <= 'h359;
    7466: romdata_int <= 'h169e;
    7467: romdata_int <= 'h40c; // Line Descriptor
    7468: romdata_int <= 'h0;
    7469: romdata_int <= 'h10ce;
    7470: romdata_int <= 'hf00;
    7471: romdata_int <= 'h40c; // Line Descriptor
    7472: romdata_int <= 'h200;
    7473: romdata_int <= 'h12fb;
    7474: romdata_int <= 'h105a;
    7475: romdata_int <= 'h40c; // Line Descriptor
    7476: romdata_int <= 'h400;
    7477: romdata_int <= 'ha3b;
    7478: romdata_int <= 'h1672;
    7479: romdata_int <= 'h40c; // Line Descriptor
    7480: romdata_int <= 'h600;
    7481: romdata_int <= 'h253;
    7482: romdata_int <= 'h745;
    7483: romdata_int <= 'h40c; // Line Descriptor
    7484: romdata_int <= 'h800;
    7485: romdata_int <= 'hec1;
    7486: romdata_int <= 'h318;
    7487: romdata_int <= 'h40c; // Line Descriptor
    7488: romdata_int <= 'ha00;
    7489: romdata_int <= 'hc5c;
    7490: romdata_int <= 'h452;
    7491: romdata_int <= 'h40c; // Line Descriptor
    7492: romdata_int <= 'hc00;
    7493: romdata_int <= 'hd3;
    7494: romdata_int <= 'h140b;
    7495: romdata_int <= 'h40c; // Line Descriptor
    7496: romdata_int <= 'he00;
    7497: romdata_int <= 'h148c;
    7498: romdata_int <= 'hac8;
    7499: romdata_int <= 'h40c; // Line Descriptor
    7500: romdata_int <= 'h1000;
    7501: romdata_int <= 'h46c;
    7502: romdata_int <= 'h129c;
    7503: romdata_int <= 'h40c; // Line Descriptor
    7504: romdata_int <= 'h1200;
    7505: romdata_int <= 'h633;
    7506: romdata_int <= 'hc0e;
    7507: romdata_int <= 'h40c; // Line Descriptor
    7508: romdata_int <= 'h1400;
    7509: romdata_int <= 'h889;
    7510: romdata_int <= 'h903;
    7511: romdata_int <= 'h50c; // Line Descriptor
    7512: romdata_int <= 'h1600;
    7513: romdata_int <= 'h1675;
    7514: romdata_int <= 'hea;
    7515: romdata_int <= 'h40a; // Line Descriptor
    7516: romdata_int <= 'ha00;
    7517: romdata_int <= 'hc59;
    7518: romdata_int <= 'ha9c;
    7519: romdata_int <= 'h40a; // Line Descriptor
    7520: romdata_int <= 'hc00;
    7521: romdata_int <= 'h6f9;
    7522: romdata_int <= 'h812;
    7523: romdata_int <= 'h40a; // Line Descriptor
    7524: romdata_int <= 'he00;
    7525: romdata_int <= 'h415;
    7526: romdata_int <= 'h141;
    7527: romdata_int <= 'h40a; // Line Descriptor
    7528: romdata_int <= 'h1000;
    7529: romdata_int <= 'he48;
    7530: romdata_int <= 'h1285;
    7531: romdata_int <= 'h40a; // Line Descriptor
    7532: romdata_int <= 'h1200;
    7533: romdata_int <= 'h1156;
    7534: romdata_int <= 'h43d;
    7535: romdata_int <= 'h40a; // Line Descriptor
    7536: romdata_int <= 'h0;
    7537: romdata_int <= 'h70a;
    7538: romdata_int <= 'hec2;
    7539: romdata_int <= 'h40a; // Line Descriptor
    7540: romdata_int <= 'h200;
    7541: romdata_int <= 'h17;
    7542: romdata_int <= 'hb0d;
    7543: romdata_int <= 'h40a; // Line Descriptor
    7544: romdata_int <= 'h400;
    7545: romdata_int <= 'haca;
    7546: romdata_int <= 'h917;
    7547: romdata_int <= 'h40a; // Line Descriptor
    7548: romdata_int <= 'h600;
    7549: romdata_int <= 'h132f;
    7550: romdata_int <= 'h61c;
    7551: romdata_int <= 'h40a; // Line Descriptor
    7552: romdata_int <= 'h800;
    7553: romdata_int <= 'h456;
    7554: romdata_int <= 'h1320;
    7555: romdata_int <= 'h40a; // Line Descriptor
    7556: romdata_int <= 'ha00;
    7557: romdata_int <= 'hc25;
    7558: romdata_int <= 'hd3;
    7559: romdata_int <= 'h40a; // Line Descriptor
    7560: romdata_int <= 'hc00;
    7561: romdata_int <= 'h8cb;
    7562: romdata_int <= 'hce4;
    7563: romdata_int <= 'h40a; // Line Descriptor
    7564: romdata_int <= 'he00;
    7565: romdata_int <= 'h25f;
    7566: romdata_int <= 'h10ce;
    7567: romdata_int <= 'h40a; // Line Descriptor
    7568: romdata_int <= 'h1000;
    7569: romdata_int <= 'h1136;
    7570: romdata_int <= 'h562;
    7571: romdata_int <= 'h40a; // Line Descriptor
    7572: romdata_int <= 'h1200;
    7573: romdata_int <= 'he1e;
    7574: romdata_int <= 'h28e;
    7575: romdata_int <= 'h40a; // Line Descriptor
    7576: romdata_int <= 'h0;
    7577: romdata_int <= 'h4e3;
    7578: romdata_int <= 'he77;
    7579: romdata_int <= 'h40a; // Line Descriptor
    7580: romdata_int <= 'h200;
    7581: romdata_int <= 'hb4;
    7582: romdata_int <= 'h148;
    7583: romdata_int <= 'h40a; // Line Descriptor
    7584: romdata_int <= 'h400;
    7585: romdata_int <= 'h221;
    7586: romdata_int <= 'h10e6;
    7587: romdata_int <= 'h40a; // Line Descriptor
    7588: romdata_int <= 'h600;
    7589: romdata_int <= 'ha2e;
    7590: romdata_int <= 'h4ff;
    7591: romdata_int <= 'h40a; // Line Descriptor
    7592: romdata_int <= 'h800;
    7593: romdata_int <= 'h1067;
    7594: romdata_int <= 'h12f7;
    7595: romdata_int <= 'h40a; // Line Descriptor
    7596: romdata_int <= 'ha00;
    7597: romdata_int <= 'h68a;
    7598: romdata_int <= 'h622;
    7599: romdata_int <= 'h40a; // Line Descriptor
    7600: romdata_int <= 'hc00;
    7601: romdata_int <= 'h809;
    7602: romdata_int <= 'hc17;
    7603: romdata_int <= 'h40a; // Line Descriptor
    7604: romdata_int <= 'he00;
    7605: romdata_int <= 'h1305;
    7606: romdata_int <= 'h20c;
    7607: romdata_int <= 'h40a; // Line Descriptor
    7608: romdata_int <= 'h1000;
    7609: romdata_int <= 'he95;
    7610: romdata_int <= 'h915;
    7611: romdata_int <= 'h40a; // Line Descriptor
    7612: romdata_int <= 'h1200;
    7613: romdata_int <= 'hcd3;
    7614: romdata_int <= 'hab9;
    7615: romdata_int <= 'h40a; // Line Descriptor
    7616: romdata_int <= 'h0;
    7617: romdata_int <= 'h448;
    7618: romdata_int <= 'h89e;
    7619: romdata_int <= 'h40a; // Line Descriptor
    7620: romdata_int <= 'h200;
    7621: romdata_int <= 'hf14;
    7622: romdata_int <= 'h2bc;
    7623: romdata_int <= 'h40a; // Line Descriptor
    7624: romdata_int <= 'h400;
    7625: romdata_int <= 'h30e;
    7626: romdata_int <= 'ha1;
    7627: romdata_int <= 'h40a; // Line Descriptor
    7628: romdata_int <= 'h600;
    7629: romdata_int <= 'h748;
    7630: romdata_int <= 'h4ad;
    7631: romdata_int <= 'h40a; // Line Descriptor
    7632: romdata_int <= 'h800;
    7633: romdata_int <= 'h1010;
    7634: romdata_int <= 'h126d;
    7635: romdata_int <= 'h40a; // Line Descriptor
    7636: romdata_int <= 'ha00;
    7637: romdata_int <= 'h933;
    7638: romdata_int <= 'h618;
    7639: romdata_int <= 'h40a; // Line Descriptor
    7640: romdata_int <= 'hc00;
    7641: romdata_int <= 'h15a;
    7642: romdata_int <= 'ha5e;
    7643: romdata_int <= 'h40a; // Line Descriptor
    7644: romdata_int <= 'he00;
    7645: romdata_int <= 'h12cc;
    7646: romdata_int <= 'hcae;
    7647: romdata_int <= 'h40a; // Line Descriptor
    7648: romdata_int <= 'h1000;
    7649: romdata_int <= 'hc38;
    7650: romdata_int <= 'he8e;
    7651: romdata_int <= 'h50a; // Line Descriptor
    7652: romdata_int <= 'h1200;
    7653: romdata_int <= 'hb62;
    7654: romdata_int <= 'h1074;
    7655: romdata_int <= 'h1808; // Line Descriptor
    7656: romdata_int <= 'h600;
    7657: romdata_int <= 'h32d;
    7658: romdata_int <= 'h63e;
    7659: romdata_int <= 'h2b9;
    7660: romdata_int <= 'h871;
    7661: romdata_int <= 'he45;
    7662: romdata_int <= 'h859;
    7663: romdata_int <= 'hc9e;
    7664: romdata_int <= 'ha29;
    7665: romdata_int <= 'h939;
    7666: romdata_int <= 'h11b;
    7667: romdata_int <= 'hcd4;
    7668: romdata_int <= 'hb5e;
    7669: romdata_int <= 'h408; // Line Descriptor
    7670: romdata_int <= 'h800;
    7671: romdata_int <= 'hf31;
    7672: romdata_int <= 'hcf0;
    7673: romdata_int <= 'h408; // Line Descriptor
    7674: romdata_int <= 'ha00;
    7675: romdata_int <= 'hc33;
    7676: romdata_int <= 'h99;
    7677: romdata_int <= 'h408; // Line Descriptor
    7678: romdata_int <= 'hc00;
    7679: romdata_int <= 'h508;
    7680: romdata_int <= 'h469;
    7681: romdata_int <= 'h408; // Line Descriptor
    7682: romdata_int <= 'he00;
    7683: romdata_int <= 'h81a;
    7684: romdata_int <= 'ha47;
    7685: romdata_int <= 'h408; // Line Descriptor
    7686: romdata_int <= 'h0;
    7687: romdata_int <= 'hf29;
    7688: romdata_int <= 'h108;
    7689: romdata_int <= 'h408; // Line Descriptor
    7690: romdata_int <= 'h200;
    7691: romdata_int <= 'hd1d;
    7692: romdata_int <= 'h925;
    7693: romdata_int <= 'h408; // Line Descriptor
    7694: romdata_int <= 'h400;
    7695: romdata_int <= 'h244;
    7696: romdata_int <= 'h666;
    7697: romdata_int <= 'h408; // Line Descriptor
    7698: romdata_int <= 'h600;
    7699: romdata_int <= 'h9e;
    7700: romdata_int <= 'he11;
    7701: romdata_int <= 'h408; // Line Descriptor
    7702: romdata_int <= 'h800;
    7703: romdata_int <= 'had4;
    7704: romdata_int <= 'h51a;
    7705: romdata_int <= 'h408; // Line Descriptor
    7706: romdata_int <= 'ha00;
    7707: romdata_int <= 'h878;
    7708: romdata_int <= 'hc14;
    7709: romdata_int <= 'h408; // Line Descriptor
    7710: romdata_int <= 'hc00;
    7711: romdata_int <= 'h40e;
    7712: romdata_int <= 'hb2d;
    7713: romdata_int <= 'h408; // Line Descriptor
    7714: romdata_int <= 'he00;
    7715: romdata_int <= 'h718;
    7716: romdata_int <= 'h20a;
    7717: romdata_int <= 'h408; // Line Descriptor
    7718: romdata_int <= 'h0;
    7719: romdata_int <= 'ha9b;
    7720: romdata_int <= 'hac5;
    7721: romdata_int <= 'h408; // Line Descriptor
    7722: romdata_int <= 'h200;
    7723: romdata_int <= 'he60;
    7724: romdata_int <= 'h215;
    7725: romdata_int <= 'h408; // Line Descriptor
    7726: romdata_int <= 'h400;
    7727: romdata_int <= 'hd4;
    7728: romdata_int <= 'h8a;
    7729: romdata_int <= 'h408; // Line Descriptor
    7730: romdata_int <= 'h600;
    7731: romdata_int <= 'h4ef;
    7732: romdata_int <= 'hf61;
    7733: romdata_int <= 'h408; // Line Descriptor
    7734: romdata_int <= 'h800;
    7735: romdata_int <= 'h842;
    7736: romdata_int <= 'h4b5;
    7737: romdata_int <= 'h408; // Line Descriptor
    7738: romdata_int <= 'ha00;
    7739: romdata_int <= 'h60b;
    7740: romdata_int <= 'hc79;
    7741: romdata_int <= 'h408; // Line Descriptor
    7742: romdata_int <= 'hc00;
    7743: romdata_int <= 'h23e;
    7744: romdata_int <= 'h916;
    7745: romdata_int <= 'h408; // Line Descriptor
    7746: romdata_int <= 'he00;
    7747: romdata_int <= 'hd22;
    7748: romdata_int <= 'h6c5;
    7749: romdata_int <= 'h408; // Line Descriptor
    7750: romdata_int <= 'h0;
    7751: romdata_int <= 'h536;
    7752: romdata_int <= 'h20;
    7753: romdata_int <= 'h408; // Line Descriptor
    7754: romdata_int <= 'h200;
    7755: romdata_int <= 'ha8b;
    7756: romdata_int <= 'ha9d;
    7757: romdata_int <= 'h408; // Line Descriptor
    7758: romdata_int <= 'h400;
    7759: romdata_int <= 'h29d;
    7760: romdata_int <= 'h4cf;
    7761: romdata_int <= 'h408; // Line Descriptor
    7762: romdata_int <= 'h600;
    7763: romdata_int <= 'hcb8;
    7764: romdata_int <= 'h299;
    7765: romdata_int <= 'h408; // Line Descriptor
    7766: romdata_int <= 'h800;
    7767: romdata_int <= 'hf39;
    7768: romdata_int <= 'h87a;
    7769: romdata_int <= 'h408; // Line Descriptor
    7770: romdata_int <= 'ha00;
    7771: romdata_int <= 'h122;
    7772: romdata_int <= 'h74e;
    7773: romdata_int <= 'h408; // Line Descriptor
    7774: romdata_int <= 'hc00;
    7775: romdata_int <= 'h636;
    7776: romdata_int <= 'hc9f;
    7777: romdata_int <= 'h408; // Line Descriptor
    7778: romdata_int <= 'he00;
    7779: romdata_int <= 'h81c;
    7780: romdata_int <= 'he3e;
    7781: romdata_int <= 'h408; // Line Descriptor
    7782: romdata_int <= 'h0;
    7783: romdata_int <= 'haeb;
    7784: romdata_int <= 'h328;
    7785: romdata_int <= 'h408; // Line Descriptor
    7786: romdata_int <= 'h200;
    7787: romdata_int <= 'h207;
    7788: romdata_int <= 'h63c;
    7789: romdata_int <= 'h408; // Line Descriptor
    7790: romdata_int <= 'h400;
    7791: romdata_int <= 'hc68;
    7792: romdata_int <= 'h483;
    7793: romdata_int <= 'h408; // Line Descriptor
    7794: romdata_int <= 'h600;
    7795: romdata_int <= 'he99;
    7796: romdata_int <= 'hcf8;
    7797: romdata_int <= 'h408; // Line Descriptor
    7798: romdata_int <= 'h800;
    7799: romdata_int <= 'h4d9;
    7800: romdata_int <= 'h808;
    7801: romdata_int <= 'h408; // Line Descriptor
    7802: romdata_int <= 'ha00;
    7803: romdata_int <= 'h12b;
    7804: romdata_int <= 'he76;
    7805: romdata_int <= 'h408; // Line Descriptor
    7806: romdata_int <= 'hc00;
    7807: romdata_int <= 'h614;
    7808: romdata_int <= 'ha50;
    7809: romdata_int <= 'h508; // Line Descriptor
    7810: romdata_int <= 'he00;
    7811: romdata_int <= 'h94a;
    7812: romdata_int <= 'hd5;
    7813: romdata_int <= 'h605; // Line Descriptor
    7814: romdata_int <= 'h0;
    7815: romdata_int <= 'h737;
    7816: romdata_int <= 'h48e;
    7817: romdata_int <= 'ha1;
    7818: romdata_int <= 'h605; // Line Descriptor
    7819: romdata_int <= 'h200;
    7820: romdata_int <= 'h122;
    7821: romdata_int <= 'h6ae;
    7822: romdata_int <= 'h50b;
    7823: romdata_int <= 'h605; // Line Descriptor
    7824: romdata_int <= 'h400;
    7825: romdata_int <= 'h35c;
    7826: romdata_int <= 'h8e1;
    7827: romdata_int <= 'h8ec;
    7828: romdata_int <= 'h605; // Line Descriptor
    7829: romdata_int <= 'h600;
    7830: romdata_int <= 'h83a;
    7831: romdata_int <= 'h2a1;
    7832: romdata_int <= 'h339;
    7833: romdata_int <= 'h605; // Line Descriptor
    7834: romdata_int <= 'h800;
    7835: romdata_int <= 'h460;
    7836: romdata_int <= 'h79;
    7837: romdata_int <= 'h6b8;
    7838: romdata_int <= 'h405; // Line Descriptor
    7839: romdata_int <= 'h0;
    7840: romdata_int <= 'h2b9;
    7841: romdata_int <= 'h73b;
    7842: romdata_int <= 'h405; // Line Descriptor
    7843: romdata_int <= 'h200;
    7844: romdata_int <= 'h49b;
    7845: romdata_int <= 'h912;
    7846: romdata_int <= 'h405; // Line Descriptor
    7847: romdata_int <= 'h400;
    7848: romdata_int <= 'h679;
    7849: romdata_int <= 'h21e;
    7850: romdata_int <= 'h405; // Line Descriptor
    7851: romdata_int <= 'h600;
    7852: romdata_int <= 'hef;
    7853: romdata_int <= 'h2a;
    7854: romdata_int <= 'h405; // Line Descriptor
    7855: romdata_int <= 'h800;
    7856: romdata_int <= 'h928;
    7857: romdata_int <= 'h48a;
    7858: romdata_int <= 'h405; // Line Descriptor
    7859: romdata_int <= 'h0;
    7860: romdata_int <= 'h455;
    7861: romdata_int <= 'h661;
    7862: romdata_int <= 'h405; // Line Descriptor
    7863: romdata_int <= 'h200;
    7864: romdata_int <= 'h6a5;
    7865: romdata_int <= 'h8e0;
    7866: romdata_int <= 'h405; // Line Descriptor
    7867: romdata_int <= 'h400;
    7868: romdata_int <= 'h8ae;
    7869: romdata_int <= 'h311;
    7870: romdata_int <= 'h405; // Line Descriptor
    7871: romdata_int <= 'h600;
    7872: romdata_int <= 'h12c;
    7873: romdata_int <= 'ha7;
    7874: romdata_int <= 'h405; // Line Descriptor
    7875: romdata_int <= 'h800;
    7876: romdata_int <= 'h32b;
    7877: romdata_int <= 'h464;
    7878: romdata_int <= 'h405; // Line Descriptor
    7879: romdata_int <= 'h0;
    7880: romdata_int <= 'h2c9;
    7881: romdata_int <= 'h354;
    7882: romdata_int <= 'h405; // Line Descriptor
    7883: romdata_int <= 'h200;
    7884: romdata_int <= 'he7;
    7885: romdata_int <= 'h413;
    7886: romdata_int <= 'h405; // Line Descriptor
    7887: romdata_int <= 'h400;
    7888: romdata_int <= 'h483;
    7889: romdata_int <= 'h718;
    7890: romdata_int <= 'h405; // Line Descriptor
    7891: romdata_int <= 'h600;
    7892: romdata_int <= 'h722;
    7893: romdata_int <= 'h87c;
    7894: romdata_int <= 'h405; // Line Descriptor
    7895: romdata_int <= 'h800;
    7896: romdata_int <= 'h855;
    7897: romdata_int <= 'h12b;
    7898: romdata_int <= 'h405; // Line Descriptor
    7899: romdata_int <= 'h0;
    7900: romdata_int <= 'h8a1;
    7901: romdata_int <= 'h4d;
    7902: romdata_int <= 'h405; // Line Descriptor
    7903: romdata_int <= 'h200;
    7904: romdata_int <= 'h449;
    7905: romdata_int <= 'h21e;
    7906: romdata_int <= 'h405; // Line Descriptor
    7907: romdata_int <= 'h400;
    7908: romdata_int <= 'h708;
    7909: romdata_int <= 'h428;
    7910: romdata_int <= 'h405; // Line Descriptor
    7911: romdata_int <= 'h600;
    7912: romdata_int <= 'hc0;
    7913: romdata_int <= 'h63f;
    7914: romdata_int <= 'h405; // Line Descriptor
    7915: romdata_int <= 'h800;
    7916: romdata_int <= 'h322;
    7917: romdata_int <= 'h8cf;
    7918: romdata_int <= 'h405; // Line Descriptor
    7919: romdata_int <= 'h0;
    7920: romdata_int <= 'h6db;
    7921: romdata_int <= 'h558;
    7922: romdata_int <= 'h405; // Line Descriptor
    7923: romdata_int <= 'h200;
    7924: romdata_int <= 'hcb;
    7925: romdata_int <= 'h71d;
    7926: romdata_int <= 'h405; // Line Descriptor
    7927: romdata_int <= 'h400;
    7928: romdata_int <= 'h2fc;
    7929: romdata_int <= 'h938;
    7930: romdata_int <= 'h405; // Line Descriptor
    7931: romdata_int <= 'h600;
    7932: romdata_int <= 'h86c;
    7933: romdata_int <= 'hee;
    7934: romdata_int <= 'h405; // Line Descriptor
    7935: romdata_int <= 'h800;
    7936: romdata_int <= 'h526;
    7937: romdata_int <= 'h2f9;
    7938: romdata_int <= 'h405; // Line Descriptor
    7939: romdata_int <= 'h0;
    7940: romdata_int <= 'h665;
    7941: romdata_int <= 'h7e;
    7942: romdata_int <= 'h405; // Line Descriptor
    7943: romdata_int <= 'h200;
    7944: romdata_int <= 'h254;
    7945: romdata_int <= 'h954;
    7946: romdata_int <= 'h405; // Line Descriptor
    7947: romdata_int <= 'h400;
    7948: romdata_int <= 'h838;
    7949: romdata_int <= 'h6b3;
    7950: romdata_int <= 'h405; // Line Descriptor
    7951: romdata_int <= 'h600;
    7952: romdata_int <= 'h44e;
    7953: romdata_int <= 'h473;
    7954: romdata_int <= 'h405; // Line Descriptor
    7955: romdata_int <= 'h800;
    7956: romdata_int <= 'he7;
    7957: romdata_int <= 'h26f;
    7958: romdata_int <= 'h405; // Line Descriptor
    7959: romdata_int <= 'h0;
    7960: romdata_int <= 'h27e;
    7961: romdata_int <= 'hc8;
    7962: romdata_int <= 'h405; // Line Descriptor
    7963: romdata_int <= 'h200;
    7964: romdata_int <= 'h492;
    7965: romdata_int <= 'h711;
    7966: romdata_int <= 'h405; // Line Descriptor
    7967: romdata_int <= 'h400;
    7968: romdata_int <= 'h709;
    7969: romdata_int <= 'h841;
    7970: romdata_int <= 'h405; // Line Descriptor
    7971: romdata_int <= 'h600;
    7972: romdata_int <= 'h12f;
    7973: romdata_int <= 'h265;
    7974: romdata_int <= 'h505; // Line Descriptor
    7975: romdata_int <= 'h800;
    7976: romdata_int <= 'h8dc;
    default: romdata_int <= 'h4ea;
  endcase
endmodule
module ldpc_edgetable(
  input        clk,
  input        rst,
  input[12:0]  romaddr,
  output[16:0] romdata
);

reg[16:0] romdata_int;

assign romdata = romdata_int;

always @( posedge rst, posedge clk )
  if( rst )
    romdata_int <= 0;
  else
  case( romaddr )
    'h0   : romdata_int = 'h10015; // Pointer for 1_4
    'h1   : romdata_int = 'h101aa; // Pointer for 1_3
    'h2   : romdata_int = 'h1038a; // Pointer for 2_5
    'h3   : romdata_int = 'h105a6; // Pointer for 1_2
    'h4   : romdata_int = 'h107c2; // Pointer for 3_5
    'h5   : romdata_int = 'h10a92; // Pointer for 2_3
    'h6   : romdata_int = 'h10cae; // Pointer for 3_4
    'h7   : romdata_int = 'h10ef7; // Pointer for 4_5
    'h8   : romdata_int = 'h1115b; // Pointer for 5_6
    'h9   : romdata_int = 'h113d1; // Pointer for 8_9
    'ha   : romdata_int = 'h115d9; // Pointer for 9_10
    'hb   : romdata_int = 'h017e3; // Pointer for 1_5s
    'hc   : romdata_int = 'h01846; // Pointer for 1_3s
    'hd   : romdata_int = 'h018be; // Pointer for 2_5s
    'he   : romdata_int = 'h01945; // Pointer for 4_9s
    'hf   : romdata_int = 'h019b3; // Pointer for 3_5s
    'h10  : romdata_int = 'h01a67; // Pointer for 2_3s
    'h11  : romdata_int = 'h01aee; // Pointer for 11_15s
    'h12  : romdata_int = 'h01b66; // Pointer for 7_9s
    'h13  : romdata_int = 'h01bd9; // Pointer for 37_45s
    'h14  : romdata_int = 'h01c5a; // Pointer for 8_9s
    'h15  : romdata_int = 'h187; // Line descriptor for 1_4
    'h16  : romdata_int = 'h4;
    'h17  : romdata_int = 'h3645;
    'h18  : romdata_int = 'h187; // Line descriptor for 1_4
    'h19  : romdata_int = 'h390b;
    'h1a  : romdata_int = 'h58f3;
    'h1b  : romdata_int = 'h187; // Line descriptor for 1_4
    'h1c  : romdata_int = 'hc0e;
    'h1d  : romdata_int = 'h1c14;
    'h1e  : romdata_int = 'h187; // Line descriptor for 1_4
    'h1f  : romdata_int = 'h1b4c;
    'h20  : romdata_int = 'h2945;
    'h21  : romdata_int = 'h187; // Line descriptor for 1_4
    'h22  : romdata_int = 'h27b;
    'h23  : romdata_int = 'h1763;
    'h24  : romdata_int = 'h187; // Line descriptor for 1_4
    'h25  : romdata_int = 'h8c9;
    'h26  : romdata_int = 'h3345;
    'h27  : romdata_int = 'h187; // Line descriptor for 1_4
    'h28  : romdata_int = 'ha67;
    'h29  : romdata_int = 'habd;
    'h2a  : romdata_int = 'h4187; // Line descriptor for 1_4
    'h2b  : romdata_int = 'h1465;
    'h2c  : romdata_int = 'h1937;
    'h2d  : romdata_int = 'h187; // Line descriptor for 1_4
    'h2e  : romdata_int = 'h311e;
    'h2f  : romdata_int = 'h46e2;
    'h30  : romdata_int = 'h187; // Line descriptor for 1_4
    'h31  : romdata_int = 'h222f;
    'h32  : romdata_int = 'h52db;
    'h33  : romdata_int = 'h187; // Line descriptor for 1_4
    'h34  : romdata_int = 'h1338;
    'h35  : romdata_int = 'h143f;
    'h36  : romdata_int = 'h187; // Line descriptor for 1_4
    'h37  : romdata_int = 'h461;
    'h38  : romdata_int = 'h183e;
    'h39  : romdata_int = 'h187; // Line descriptor for 1_4
    'h3a  : romdata_int = 'h10df;
    'h3b  : romdata_int = 'h1ea4;
    'h3c  : romdata_int = 'h187; // Line descriptor for 1_4
    'h3d  : romdata_int = 'h1ced;
    'h3e  : romdata_int = 'h54f3;
    'h3f  : romdata_int = 'h4187; // Line descriptor for 1_4
    'h40  : romdata_int = 'h1690;
    'h41  : romdata_int = 'h3a36;
    'h42  : romdata_int = 'h187; // Line descriptor for 1_4
    'h43  : romdata_int = 'h89;
    'h44  : romdata_int = 'h4e0;
    'h45  : romdata_int = 'h187; // Line descriptor for 1_4
    'h46  : romdata_int = 'h2e;
    'h47  : romdata_int = 'hf48;
    'h48  : romdata_int = 'h187; // Line descriptor for 1_4
    'h49  : romdata_int = 'h1144;
    'h4a  : romdata_int = 'h185c;
    'h4b  : romdata_int = 'h187; // Line descriptor for 1_4
    'h4c  : romdata_int = 'h12ce;
    'h4d  : romdata_int = 'h507e;
    'h4e  : romdata_int = 'h187; // Line descriptor for 1_4
    'h4f  : romdata_int = 'h1135;
    'h50  : romdata_int = 'h18c3;
    'h51  : romdata_int = 'h187; // Line descriptor for 1_4
    'h52  : romdata_int = 'h1746;
    'h53  : romdata_int = 'h3c60;
    'h54  : romdata_int = 'h4187; // Line descriptor for 1_4
    'h55  : romdata_int = 'h1ccb;
    'h56  : romdata_int = 'h2eb3;
    'h57  : romdata_int = 'h187; // Line descriptor for 1_4
    'h58  : romdata_int = 'h2b9;
    'h59  : romdata_int = 'h4711;
    'h5a  : romdata_int = 'h187; // Line descriptor for 1_4
    'h5b  : romdata_int = 'h14c0;
    'h5c  : romdata_int = 'h4838;
    'h5d  : romdata_int = 'h187; // Line descriptor for 1_4
    'h5e  : romdata_int = 'hd4d;
    'h5f  : romdata_int = 'h10d6;
    'h60  : romdata_int = 'h187; // Line descriptor for 1_4
    'h61  : romdata_int = 'haa6;
    'h62  : romdata_int = 'h1b15;
    'h63  : romdata_int = 'h187; // Line descriptor for 1_4
    'h64  : romdata_int = 'h2303;
    'h65  : romdata_int = 'h44b5;
    'h66  : romdata_int = 'h187; // Line descriptor for 1_4
    'h67  : romdata_int = 'h642;
    'h68  : romdata_int = 'h8d5;
    'h69  : romdata_int = 'h4187; // Line descriptor for 1_4
    'h6a  : romdata_int = 'hf2a;
    'h6b  : romdata_int = 'h1d1f;
    'h6c  : romdata_int = 'h187; // Line descriptor for 1_4
    'h6d  : romdata_int = 'h137;
    'h6e  : romdata_int = 'h46b;
    'h6f  : romdata_int = 'h187; // Line descriptor for 1_4
    'h70  : romdata_int = 'hd38;
    'h71  : romdata_int = 'h3c7d;
    'h72  : romdata_int = 'h187; // Line descriptor for 1_4
    'h73  : romdata_int = 'h84a;
    'h74  : romdata_int = 'haf2;
    'h75  : romdata_int = 'h187; // Line descriptor for 1_4
    'h76  : romdata_int = 'h30e5;
    'h77  : romdata_int = 'h48b4;
    'h78  : romdata_int = 'h187; // Line descriptor for 1_4
    'h79  : romdata_int = 'h16b4;
    'h7a  : romdata_int = 'h3307;
    'h7b  : romdata_int = 'h187; // Line descriptor for 1_4
    'h7c  : romdata_int = 'h312;
    'h7d  : romdata_int = 'h10a0;
    'h7e  : romdata_int = 'h4187; // Line descriptor for 1_4
    'h7f  : romdata_int = 'h14e5;
    'h80  : romdata_int = 'h5045;
    'h81  : romdata_int = 'h187; // Line descriptor for 1_4
    'h82  : romdata_int = 'h92b;
    'h83  : romdata_int = 'hcab;
    'h84  : romdata_int = 'h187; // Line descriptor for 1_4
    'h85  : romdata_int = 'h12fd;
    'h86  : romdata_int = 'h299;
    'h87  : romdata_int = 'h187; // Line descriptor for 1_4
    'h88  : romdata_int = 'h728;
    'h89  : romdata_int = 'h36a2;
    'h8a  : romdata_int = 'h187; // Line descriptor for 1_4
    'h8b  : romdata_int = 'h1221;
    'h8c  : romdata_int = 'h266a;
    'h8d  : romdata_int = 'h187; // Line descriptor for 1_4
    'h8e  : romdata_int = 'hb2c;
    'h8f  : romdata_int = 'h4241;
    'h90  : romdata_int = 'h187; // Line descriptor for 1_4
    'h91  : romdata_int = 'h1a64;
    'h92  : romdata_int = 'h1aad;
    'h93  : romdata_int = 'h4187; // Line descriptor for 1_4
    'h94  : romdata_int = 'hb0;
    'h95  : romdata_int = 'h208f;
    'h96  : romdata_int = 'h187; // Line descriptor for 1_4
    'h97  : romdata_int = 'h2a3f;
    'h98  : romdata_int = 'h4a03;
    'h99  : romdata_int = 'h187; // Line descriptor for 1_4
    'h9a  : romdata_int = 'h455;
    'h9b  : romdata_int = 'h121c;
    'h9c  : romdata_int = 'h187; // Line descriptor for 1_4
    'h9d  : romdata_int = 'ha88;
    'h9e  : romdata_int = 'h109b;
    'h9f  : romdata_int = 'h187; // Line descriptor for 1_4
    'ha0  : romdata_int = 'hc25;
    'ha1  : romdata_int = 'h18ca;
    'ha2  : romdata_int = 'h187; // Line descriptor for 1_4
    'ha3  : romdata_int = 'he66;
    'ha4  : romdata_int = 'h2767;
    'ha5  : romdata_int = 'h187; // Line descriptor for 1_4
    'ha6  : romdata_int = 'h167e;
    'ha7  : romdata_int = 'hc4c;
    'ha8  : romdata_int = 'h4187; // Line descriptor for 1_4
    'ha9  : romdata_int = 'h168f;
    'haa  : romdata_int = 'h1b58;
    'hab  : romdata_int = 'h187; // Line descriptor for 1_4
    'hac  : romdata_int = 'h864;
    'had  : romdata_int = 'h3ea6;
    'hae  : romdata_int = 'h187; // Line descriptor for 1_4
    'haf  : romdata_int = 'hf16;
    'hb0  : romdata_int = 'h1a17;
    'hb1  : romdata_int = 'h187; // Line descriptor for 1_4
    'hb2  : romdata_int = 'h936;
    'hb3  : romdata_int = 'h1054;
    'hb4  : romdata_int = 'h187; // Line descriptor for 1_4
    'hb5  : romdata_int = 'h10b;
    'hb6  : romdata_int = 'h1b06;
    'hb7  : romdata_int = 'h187; // Line descriptor for 1_4
    'hb8  : romdata_int = 'h1670;
    'hb9  : romdata_int = 'h2e97;
    'hba  : romdata_int = 'h187; // Line descriptor for 1_4
    'hbb  : romdata_int = 'h2cb1;
    'hbc  : romdata_int = 'h4e6;
    'hbd  : romdata_int = 'h4187; // Line descriptor for 1_4
    'hbe  : romdata_int = 'h2cd5;
    'hbf  : romdata_int = 'h4ac8;
    'hc0  : romdata_int = 'h187; // Line descriptor for 1_4
    'hc1  : romdata_int = 'hc41;
    'hc2  : romdata_int = 'h1319;
    'hc3  : romdata_int = 'h187; // Line descriptor for 1_4
    'hc4  : romdata_int = 'h86;
    'hc5  : romdata_int = 'h4ce8;
    'hc6  : romdata_int = 'h187; // Line descriptor for 1_4
    'hc7  : romdata_int = 'h51e;
    'hc8  : romdata_int = 'h62d;
    'hc9  : romdata_int = 'h187; // Line descriptor for 1_4
    'hca  : romdata_int = 'h8;
    'hcb  : romdata_int = 'he58;
    'hcc  : romdata_int = 'h187; // Line descriptor for 1_4
    'hcd  : romdata_int = 'h161f;
    'hce  : romdata_int = 'h4e10;
    'hcf  : romdata_int = 'h187; // Line descriptor for 1_4
    'hd0  : romdata_int = 'h33b;
    'hd1  : romdata_int = 'h1e3d;
    'hd2  : romdata_int = 'h4187; // Line descriptor for 1_4
    'hd3  : romdata_int = 'h1d3d;
    'hd4  : romdata_int = 'h5280;
    'hd5  : romdata_int = 'h187; // Line descriptor for 1_4
    'hd6  : romdata_int = 'h1a42;
    'hd7  : romdata_int = 'h72c;
    'hd8  : romdata_int = 'h187; // Line descriptor for 1_4
    'hd9  : romdata_int = 'hc75;
    'hda  : romdata_int = 'h173f;
    'hdb  : romdata_int = 'h187; // Line descriptor for 1_4
    'hdc  : romdata_int = 'h1a2b;
    'hdd  : romdata_int = 'h435e;
    'hde  : romdata_int = 'h187; // Line descriptor for 1_4
    'hdf  : romdata_int = 'h1030;
    'he0  : romdata_int = 'h1887;
    'he1  : romdata_int = 'h187; // Line descriptor for 1_4
    'he2  : romdata_int = 'h1623;
    'he3  : romdata_int = 'h4c59;
    'he4  : romdata_int = 'h187; // Line descriptor for 1_4
    'he5  : romdata_int = 'h122a;
    'he6  : romdata_int = 'h4606;
    'he7  : romdata_int = 'h4187; // Line descriptor for 1_4
    'he8  : romdata_int = 'h10d0;
    'he9  : romdata_int = 'h4ca0;
    'hea  : romdata_int = 'h187; // Line descriptor for 1_4
    'heb  : romdata_int = 'h4d5;
    'hec  : romdata_int = 'h3434;
    'hed  : romdata_int = 'h187; // Line descriptor for 1_4
    'hee  : romdata_int = 'h83b;
    'hef  : romdata_int = 'h446f;
    'hf0  : romdata_int = 'h187; // Line descriptor for 1_4
    'hf1  : romdata_int = 'hb22;
    'hf2  : romdata_int = 'he4d;
    'hf3  : romdata_int = 'h187; // Line descriptor for 1_4
    'hf4  : romdata_int = 'h48a;
    'hf5  : romdata_int = 'h862;
    'hf6  : romdata_int = 'h187; // Line descriptor for 1_4
    'hf7  : romdata_int = 'h12c9;
    'hf8  : romdata_int = 'h1522;
    'hf9  : romdata_int = 'h187; // Line descriptor for 1_4
    'hfa  : romdata_int = 'h1958;
    'hfb  : romdata_int = 'h4e85;
    'hfc  : romdata_int = 'h4187; // Line descriptor for 1_4
    'hfd  : romdata_int = 'h18db;
    'hfe  : romdata_int = 'ha5c;
    'hff  : romdata_int = 'h187; // Line descriptor for 1_4
    'h100 : romdata_int = 'h1d1d;
    'h101 : romdata_int = 'h346f;
    'h102 : romdata_int = 'h187; // Line descriptor for 1_4
    'h103 : romdata_int = 'h168c;
    'h104 : romdata_int = 'h4e08;
    'h105 : romdata_int = 'h187; // Line descriptor for 1_4
    'h106 : romdata_int = 'h954;
    'h107 : romdata_int = 'hd52;
    'h108 : romdata_int = 'h187; // Line descriptor for 1_4
    'h109 : romdata_int = 'h16da;
    'h10a : romdata_int = 'h22f8;
    'h10b : romdata_int = 'h187; // Line descriptor for 1_4
    'h10c : romdata_int = 'h24dc;
    'h10d : romdata_int = 'h4049;
    'h10e : romdata_int = 'h187; // Line descriptor for 1_4
    'h10f : romdata_int = 'h673;
    'h110 : romdata_int = 'hb49;
    'h111 : romdata_int = 'h4187; // Line descriptor for 1_4
    'h112 : romdata_int = 'h279;
    'h113 : romdata_int = 'h3eaf;
    'h114 : romdata_int = 'h187; // Line descriptor for 1_4
    'h115 : romdata_int = 'h1006;
    'h116 : romdata_int = 'h4149;
    'h117 : romdata_int = 'h187; // Line descriptor for 1_4
    'h118 : romdata_int = 'h890;
    'h119 : romdata_int = 'h10be;
    'h11a : romdata_int = 'h187; // Line descriptor for 1_4
    'h11b : romdata_int = 'hef3;
    'h11c : romdata_int = 'h303c;
    'h11d : romdata_int = 'h187; // Line descriptor for 1_4
    'h11e : romdata_int = 'h2b8;
    'h11f : romdata_int = 'h4a5;
    'h120 : romdata_int = 'h187; // Line descriptor for 1_4
    'h121 : romdata_int = 'h187b;
    'h122 : romdata_int = 'h9a;
    'h123 : romdata_int = 'h187; // Line descriptor for 1_4
    'h124 : romdata_int = 'h1031;
    'h125 : romdata_int = 'h1845;
    'h126 : romdata_int = 'h4187; // Line descriptor for 1_4
    'h127 : romdata_int = 'h302;
    'h128 : romdata_int = 'h3857;
    'h129 : romdata_int = 'h187; // Line descriptor for 1_4
    'h12a : romdata_int = 'h3b26;
    'h12b : romdata_int = 'h4a22;
    'h12c : romdata_int = 'h187; // Line descriptor for 1_4
    'h12d : romdata_int = 'h24da;
    'h12e : romdata_int = 'h5555;
    'h12f : romdata_int = 'h187; // Line descriptor for 1_4
    'h130 : romdata_int = 'h18ee;
    'h131 : romdata_int = 'h6e5;
    'h132 : romdata_int = 'h187; // Line descriptor for 1_4
    'h133 : romdata_int = 'h24e4;
    'h134 : romdata_int = 'h52b5;
    'h135 : romdata_int = 'h187; // Line descriptor for 1_4
    'h136 : romdata_int = 'h1906;
    'h137 : romdata_int = 'h1eb3;
    'h138 : romdata_int = 'h187; // Line descriptor for 1_4
    'h139 : romdata_int = 'h1c9a;
    'h13a : romdata_int = 'h2af5;
    'h13b : romdata_int = 'h4187; // Line descriptor for 1_4
    'h13c : romdata_int = 'hf58;
    'h13d : romdata_int = 'h2644;
    'h13e : romdata_int = 'h187; // Line descriptor for 1_4
    'h13f : romdata_int = 'h467;
    'h140 : romdata_int = 'h1308;
    'h141 : romdata_int = 'h187; // Line descriptor for 1_4
    'h142 : romdata_int = 'h6a7;
    'h143 : romdata_int = 'h1418;
    'h144 : romdata_int = 'h187; // Line descriptor for 1_4
    'h145 : romdata_int = 'he1a;
    'h146 : romdata_int = 'h3e52;
    'h147 : romdata_int = 'h187; // Line descriptor for 1_4
    'h148 : romdata_int = 'h1a35;
    'h149 : romdata_int = 'h5898;
    'h14a : romdata_int = 'h187; // Line descriptor for 1_4
    'h14b : romdata_int = 'h27f;
    'h14c : romdata_int = 'h14eb;
    'h14d : romdata_int = 'h187; // Line descriptor for 1_4
    'h14e : romdata_int = 'hd5;
    'h14f : romdata_int = 'hb27;
    'h150 : romdata_int = 'h4187; // Line descriptor for 1_4
    'h151 : romdata_int = 'h3628;
    'h152 : romdata_int = 'h511e;
    'h153 : romdata_int = 'h187; // Line descriptor for 1_4
    'h154 : romdata_int = 'h14fd;
    'h155 : romdata_int = 'h3af9;
    'h156 : romdata_int = 'h187; // Line descriptor for 1_4
    'h157 : romdata_int = 'h1d31;
    'h158 : romdata_int = 'h1440;
    'h159 : romdata_int = 'h187; // Line descriptor for 1_4
    'h15a : romdata_int = 'h15c;
    'h15b : romdata_int = 'hd4f;
    'h15c : romdata_int = 'h187; // Line descriptor for 1_4
    'h15d : romdata_int = 'h8b6;
    'h15e : romdata_int = 'h38f3;
    'h15f : romdata_int = 'h187; // Line descriptor for 1_4
    'h160 : romdata_int = 'h1cc4;
    'h161 : romdata_int = 'h5959;
    'h162 : romdata_int = 'h187; // Line descriptor for 1_4
    'h163 : romdata_int = 'hc8f;
    'h164 : romdata_int = 'h1408;
    'h165 : romdata_int = 'h4187; // Line descriptor for 1_4
    'h166 : romdata_int = 'h2e1d;
    'h167 : romdata_int = 'h5711;
    'h168 : romdata_int = 'h187; // Line descriptor for 1_4
    'h169 : romdata_int = 'h1233;
    'h16a : romdata_int = 'hc70;
    'h16b : romdata_int = 'h187; // Line descriptor for 1_4
    'h16c : romdata_int = 'h67c;
    'h16d : romdata_int = 'h6a4;
    'h16e : romdata_int = 'h187; // Line descriptor for 1_4
    'h16f : romdata_int = 'h1250;
    'h170 : romdata_int = 'h281e;
    'h171 : romdata_int = 'h187; // Line descriptor for 1_4
    'h172 : romdata_int = 'hae;
    'h173 : romdata_int = 'h40ff;
    'h174 : romdata_int = 'h187; // Line descriptor for 1_4
    'h175 : romdata_int = 'h29b;
    'h176 : romdata_int = 'h1a73;
    'h177 : romdata_int = 'h187; // Line descriptor for 1_4
    'h178 : romdata_int = 'h27c;
    'h179 : romdata_int = 'h145d;
    'h17a : romdata_int = 'h4187; // Line descriptor for 1_4
    'h17b : romdata_int = 'h40d;
    'h17c : romdata_int = 'h1c0a;
    'h17d : romdata_int = 'h187; // Line descriptor for 1_4
    'h17e : romdata_int = 'h2afe;
    'h17f : romdata_int = 'h5687;
    'h180 : romdata_int = 'h187; // Line descriptor for 1_4
    'h181 : romdata_int = 'h147b;
    'h182 : romdata_int = 'h3551;
    'h183 : romdata_int = 'h187; // Line descriptor for 1_4
    'h184 : romdata_int = 'h6a6;
    'h185 : romdata_int = 'h4550;
    'h186 : romdata_int = 'h187; // Line descriptor for 1_4
    'h187 : romdata_int = 'h2049;
    'h188 : romdata_int = 'h5696;
    'h189 : romdata_int = 'h187; // Line descriptor for 1_4
    'h18a : romdata_int = 'heee;
    'h18b : romdata_int = 'h54e5;
    'h18c : romdata_int = 'h187; // Line descriptor for 1_4
    'h18d : romdata_int = 'h1cc9;
    'h18e : romdata_int = 'h2ca6;
    'h18f : romdata_int = 'h4187; // Line descriptor for 1_4
    'h190 : romdata_int = 'h8f2;
    'h191 : romdata_int = 'h2919;
    'h192 : romdata_int = 'h187; // Line descriptor for 1_4
    'h193 : romdata_int = 'h20cd;
    'h194 : romdata_int = 'h3cdd;
    'h195 : romdata_int = 'h187; // Line descriptor for 1_4
    'h196 : romdata_int = 'hb01;
    'h197 : romdata_int = 'h1ac5;
    'h198 : romdata_int = 'h187; // Line descriptor for 1_4
    'h199 : romdata_int = 'h1d5b;
    'h19a : romdata_int = 'h329e;
    'h19b : romdata_int = 'h187; // Line descriptor for 1_4
    'h19c : romdata_int = 'he0a;
    'h19d : romdata_int = 'h4267;
    'h19e : romdata_int = 'h187; // Line descriptor for 1_4
    'h19f : romdata_int = 'h643;
    'h1a0 : romdata_int = 'ha48;
    'h1a1 : romdata_int = 'h187; // Line descriptor for 1_4
    'h1a2 : romdata_int = 'h6b0;
    'h1a3 : romdata_int = 'h12a2;
    'h1a4 : romdata_int = 'h4187; // Line descriptor for 1_4
    'h1a5 : romdata_int = 'h238;
    'h1a6 : romdata_int = 'he32;
    'h1a7 : romdata_int = 'h2187; // Line descriptor for 1_4
    'h1a8 : romdata_int = 'h528;
    'h1a9 : romdata_int = 'h4862;
    'h1aa : romdata_int = 'h278; // Line descriptor for 1_3
    'h1ab : romdata_int = 'h2e;
    'h1ac : romdata_int = 'hb0;
    'h1ad : romdata_int = 'h5939;
    'h1ae : romdata_int = 'h278; // Line descriptor for 1_3
    'h1af : romdata_int = 'h46e4;
    'h1b0 : romdata_int = 'h5cb8;
    'h1b1 : romdata_int = 'h6cec;
    'h1b2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h1b3 : romdata_int = 'hc8f;
    'h1b4 : romdata_int = 'h20f3;
    'h1b5 : romdata_int = 'h371c;
    'h1b6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h1b7 : romdata_int = 'h27b;
    'h1b8 : romdata_int = 'h194c;
    'h1b9 : romdata_int = 'h5cd1;
    'h1ba : romdata_int = 'h4278; // Line descriptor for 1_3
    'h1bb : romdata_int = 'h1563;
    'h1bc : romdata_int = 'h1a14;
    'h1bd : romdata_int = 'h2f59;
    'h1be : romdata_int = 'h278; // Line descriptor for 1_3
    'h1bf : romdata_int = 'h8c9;
    'h1c0 : romdata_int = 'h2256;
    'h1c1 : romdata_int = 'h2410;
    'h1c2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h1c3 : romdata_int = 'ha67;
    'h1c4 : romdata_int = 'habd;
    'h1c5 : romdata_int = 'h1f07;
    'h1c6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h1c7 : romdata_int = 'h1265;
    'h1c8 : romdata_int = 'h2480;
    'h1c9 : romdata_int = 'h5e43;
    'h1ca : romdata_int = 'h278; // Line descriptor for 1_3
    'h1cb : romdata_int = 'h2a91;
    'h1cc : romdata_int = 'h2c85;
    'h1cd : romdata_int = 'h454a;
    'h1ce : romdata_int = 'h4278; // Line descriptor for 1_3
    'h1cf : romdata_int = 'h1321;
    'h1d0 : romdata_int = 'h2036;
    'h1d1 : romdata_int = 'h2ee3;
    'h1d2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h1d3 : romdata_int = 'h461;
    'h1d4 : romdata_int = 'h26b1;
    'h1d5 : romdata_int = 'h5b07;
    'h1d6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h1d7 : romdata_int = 'h206c;
    'h1d8 : romdata_int = 'h1138;
    'h1d9 : romdata_int = 'h123f;
    'h1da : romdata_int = 'h278; // Line descriptor for 1_3
    'h1db : romdata_int = 'h1c97;
    'h1dc : romdata_int = 'h6c29;
    'h1dd : romdata_int = 'h2137;
    'h1de : romdata_int = 'h278; // Line descriptor for 1_3
    'h1df : romdata_int = 'h86;
    'h1e0 : romdata_int = 'h163e;
    'h1e1 : romdata_int = 'h1490;
    'h1e2 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h1e3 : romdata_int = 'h2d43;
    'h1e4 : romdata_int = 'h4e0;
    'h1e5 : romdata_int = 'h89;
    'h1e6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h1e7 : romdata_int = 'hf48;
    'h1e8 : romdata_int = 'h165c;
    'h1e9 : romdata_int = 'h5877;
    'h1ea : romdata_int = 'h278; // Line descriptor for 1_3
    'h1eb : romdata_int = 'h2206;
    'h1ec : romdata_int = 'h680a;
    'h1ed : romdata_int = 'h7242;
    'h1ee : romdata_int = 'h278; // Line descriptor for 1_3
    'h1ef : romdata_int = 'h1aed;
    'h1f0 : romdata_int = 'h44b0;
    'h1f1 : romdata_int = 'h46f5;
    'h1f2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h1f3 : romdata_int = 'hf05;
    'h1f4 : romdata_int = 'h10ce;
    'h1f5 : romdata_int = 'h7458;
    'h1f6 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h1f7 : romdata_int = 'h1546;
    'h1f8 : romdata_int = 'h2ced;
    'h1f9 : romdata_int = 'h5cd3;
    'h1fa : romdata_int = 'h278; // Line descriptor for 1_3
    'h1fb : romdata_int = 'h1c3f;
    'h1fc : romdata_int = 'h414c;
    'h1fd : romdata_int = 'h1461;
    'h1fe : romdata_int = 'h278; // Line descriptor for 1_3
    'h1ff : romdata_int = 'hb53;
    'h200 : romdata_int = 'h16c3;
    'h201 : romdata_int = 'h20ee;
    'h202 : romdata_int = 'h278; // Line descriptor for 1_3
    'h203 : romdata_int = 'h2b9;
    'h204 : romdata_int = 'hea1;
    'h205 : romdata_int = 'h1915;
    'h206 : romdata_int = 'h278; // Line descriptor for 1_3
    'h207 : romdata_int = 'h642;
    'h208 : romdata_int = 'h2249;
    'h209 : romdata_int = 'h3a94;
    'h20a : romdata_int = 'h4278; // Line descriptor for 1_3
    'h20b : romdata_int = 'h12c0;
    'h20c : romdata_int = 'h4aa0;
    'h20d : romdata_int = 'h569b;
    'h20e : romdata_int = 'h278; // Line descriptor for 1_3
    'h20f : romdata_int = 'hc25;
    'h210 : romdata_int = 'h1e9e;
    'h211 : romdata_int = 'h24ee;
    'h212 : romdata_int = 'h278; // Line descriptor for 1_3
    'h213 : romdata_int = 'h4;
    'h214 : romdata_int = 'haa6;
    'h215 : romdata_int = 'h10fe;
    'h216 : romdata_int = 'h278; // Line descriptor for 1_3
    'h217 : romdata_int = 'h46b;
    'h218 : romdata_int = 'hf2a;
    'h219 : romdata_int = 'h6e22;
    'h21a : romdata_int = 'h278; // Line descriptor for 1_3
    'h21b : romdata_int = 'h8d5;
    'h21c : romdata_int = 'h2260;
    'h21d : romdata_int = 'h7343;
    'h21e : romdata_int = 'h4278; // Line descriptor for 1_3
    'h21f : romdata_int = 'h1abb;
    'h220 : romdata_int = 'h28eb;
    'h221 : romdata_int = 'h52d6;
    'h222 : romdata_int = 'h278; // Line descriptor for 1_3
    'h223 : romdata_int = 'h312;
    'h224 : romdata_int = 'hd52;
    'h225 : romdata_int = 'h2091;
    'h226 : romdata_int = 'h278; // Line descriptor for 1_3
    'h227 : romdata_int = 'h92b;
    'h228 : romdata_int = 'h1b1f;
    'h229 : romdata_int = 'h774b;
    'h22a : romdata_int = 'h278; // Line descriptor for 1_3
    'h22b : romdata_int = 'haf2;
    'h22c : romdata_int = 'hc0e;
    'h22d : romdata_int = 'h273b;
    'h22e : romdata_int = 'h278; // Line descriptor for 1_3
    'h22f : romdata_int = 'h4205;
    'h230 : romdata_int = 'h608e;
    'h231 : romdata_int = 'h76d3;
    'h232 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h233 : romdata_int = 'h728;
    'h234 : romdata_int = 'h3167;
    'h235 : romdata_int = 'h6b66;
    'h236 : romdata_int = 'h278; // Line descriptor for 1_3
    'h237 : romdata_int = 'hb2c;
    'h238 : romdata_int = 'h1e39;
    'h239 : romdata_int = 'h1e8b;
    'h23a : romdata_int = 'h278; // Line descriptor for 1_3
    'h23b : romdata_int = 'h247e;
    'h23c : romdata_int = 'h5162;
    'h23d : romdata_int = 'h68d2;
    'h23e : romdata_int = 'h278; // Line descriptor for 1_3
    'h23f : romdata_int = 'h101c;
    'h240 : romdata_int = 'h10fd;
    'h241 : romdata_int = 'h3274;
    'h242 : romdata_int = 'h278; // Line descriptor for 1_3
    'h243 : romdata_int = 'h9a;
    'h244 : romdata_int = 'hd4f;
    'h245 : romdata_int = 'h12e5;
    'h246 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h247 : romdata_int = 'h16ca;
    'h248 : romdata_int = 'h1cfc;
    'h249 : romdata_int = 'h1cfe;
    'h24a : romdata_int = 'h278; // Line descriptor for 1_3
    'h24b : romdata_int = 'h147e;
    'h24c : romdata_int = 'h18ad;
    'h24d : romdata_int = 'h2430;
    'h24e : romdata_int = 'h278; // Line descriptor for 1_3
    'h24f : romdata_int = 'h455;
    'h250 : romdata_int = 'h200e;
    'h251 : romdata_int = 'h6a48;
    'h252 : romdata_int = 'h278; // Line descriptor for 1_3
    'h253 : romdata_int = 'he66;
    'h254 : romdata_int = 'h2458;
    'h255 : romdata_int = 'h7622;
    'h256 : romdata_int = 'h278; // Line descriptor for 1_3
    'h257 : romdata_int = 'h864;
    'h258 : romdata_int = 'h1817;
    'h259 : romdata_int = 'h1d38;
    'h25a : romdata_int = 'h4278; // Line descriptor for 1_3
    'h25b : romdata_int = 'h24b5;
    'h25c : romdata_int = 'h3d4c;
    'h25d : romdata_int = 'h6052;
    'h25e : romdata_int = 'h278; // Line descriptor for 1_3
    'h25f : romdata_int = 'ha88;
    'h260 : romdata_int = 'h160b;
    'h261 : romdata_int = 'h5887;
    'h262 : romdata_int = 'h278; // Line descriptor for 1_3
    'h263 : romdata_int = 'h1470;
    'h264 : romdata_int = 'h1ee5;
    'h265 : romdata_int = 'h4e13;
    'h266 : romdata_int = 'h278; // Line descriptor for 1_3
    'h267 : romdata_int = 'hae;
    'h268 : romdata_int = 'h2238;
    'h269 : romdata_int = 'h647b;
    'h26a : romdata_int = 'h278; // Line descriptor for 1_3
    'h26b : romdata_int = 'h1958;
    'h26c : romdata_int = 'h24a8;
    'h26d : romdata_int = 'h7424;
    'h26e : romdata_int = 'h4278; // Line descriptor for 1_3
    'h26f : romdata_int = 'h491;
    'h270 : romdata_int = 'hf16;
    'h271 : romdata_int = 'h6d1d;
    'h272 : romdata_int = 'h278; // Line descriptor for 1_3
    'h273 : romdata_int = 'h2057;
    'h274 : romdata_int = 'h1842;
    'h275 : romdata_int = 'h2465;
    'h276 : romdata_int = 'h278; // Line descriptor for 1_3
    'h277 : romdata_int = 'hd5;
    'h278 : romdata_int = 'h1b3d;
    'h279 : romdata_int = 'h20f4;
    'h27a : romdata_int = 'h278; // Line descriptor for 1_3
    'h27b : romdata_int = 'h51e;
    'h27c : romdata_int = 'h1e3c;
    'h27d : romdata_int = 'h3633;
    'h27e : romdata_int = 'h278; // Line descriptor for 1_3
    'h27f : romdata_int = 'h10b;
    'h280 : romdata_int = 'h936;
    'h281 : romdata_int = 'h26d4;
    'h282 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h283 : romdata_int = 'h3a54;
    'h284 : romdata_int = 'h4af2;
    'h285 : romdata_int = 'h6486;
    'h286 : romdata_int = 'h278; // Line descriptor for 1_3
    'h287 : romdata_int = 'h1119;
    'h288 : romdata_int = 'h1687;
    'h289 : romdata_int = 'h182b;
    'h28a : romdata_int = 'h278; // Line descriptor for 1_3
    'h28b : romdata_int = 'h72c;
    'h28c : romdata_int = 'h33b;
    'h28d : romdata_int = 'h5747;
    'h28e : romdata_int = 'h278; // Line descriptor for 1_3
    'h28f : romdata_int = 'hcab;
    'h290 : romdata_int = 'h1706;
    'h291 : romdata_int = 'h62d;
    'h292 : romdata_int = 'h278; // Line descriptor for 1_3
    'h293 : romdata_int = 'h141f;
    'h294 : romdata_int = 'h22d8;
    'h295 : romdata_int = 'h649b;
    'h296 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h297 : romdata_int = 'h28cf;
    'h298 : romdata_int = 'h3229;
    'h299 : romdata_int = 'h4818;
    'h29a : romdata_int = 'h278; // Line descriptor for 1_3
    'h29b : romdata_int = 'h1f66;
    'h29c : romdata_int = 'h1f4d;
    'h29d : romdata_int = 'h102a;
    'h29e : romdata_int = 'h278; // Line descriptor for 1_3
    'h29f : romdata_int = 'h1e81;
    'h2a0 : romdata_int = 'h391c;
    'h2a1 : romdata_int = 'he4d;
    'h2a2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2a3 : romdata_int = 'h4d5;
    'h2a4 : romdata_int = 'h223a;
    'h2a5 : romdata_int = 'h6ace;
    'h2a6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2a7 : romdata_int = 'h83b;
    'h2a8 : romdata_int = 'hb22;
    'h2a9 : romdata_int = 'h153f;
    'h2aa : romdata_int = 'h4278; // Line descriptor for 1_3
    'h2ab : romdata_int = 'h48a;
    'h2ac : romdata_int = 'h4e70;
    'h2ad : romdata_int = 'h6712;
    'h2ae : romdata_int = 'h278; // Line descriptor for 1_3
    'h2af : romdata_int = 'h1423;
    'h2b0 : romdata_int = 'h2ee4;
    'h2b1 : romdata_int = 'h3a7a;
    'h2b2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2b3 : romdata_int = 'ha5c;
    'h2b4 : romdata_int = 'h1758;
    'h2b5 : romdata_int = 'h1f1e;
    'h2b6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2b7 : romdata_int = 'h862;
    'h2b8 : romdata_int = 'h148c;
    'h2b9 : romdata_int = 'h26f3;
    'h2ba : romdata_int = 'h278; // Line descriptor for 1_3
    'h2bb : romdata_int = 'h10c9;
    'h2bc : romdata_int = 'h167b;
    'h2bd : romdata_int = 'h7078;
    'h2be : romdata_int = 'h4278; // Line descriptor for 1_3
    'h2bf : romdata_int = 'h14da;
    'h2c0 : romdata_int = 'h1f45;
    'h2c1 : romdata_int = 'h3157;
    'h2c2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2c3 : romdata_int = 'h954;
    'h2c4 : romdata_int = 'h16db;
    'h2c5 : romdata_int = 'h1d45;
    'h2c6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2c7 : romdata_int = 'h2203;
    'h2c8 : romdata_int = 'h2445;
    'h2c9 : romdata_int = 'h40f2;
    'h2ca : romdata_int = 'h278; // Line descriptor for 1_3
    'h2cb : romdata_int = 'h852;
    'h2cc : romdata_int = 'h3523;
    'h2cd : romdata_int = 'h4317;
    'h2ce : romdata_int = 'h278; // Line descriptor for 1_3
    'h2cf : romdata_int = 'h673;
    'h2d0 : romdata_int = 'h1c1e;
    'h2d1 : romdata_int = 'h246e;
    'h2d2 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h2d3 : romdata_int = 'h279;
    'h2d4 : romdata_int = 'hd4d;
    'h2d5 : romdata_int = 'h1645;
    'h2d6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2d7 : romdata_int = 'h6f3;
    'h2d8 : romdata_int = 'h22b4;
    'h2d9 : romdata_int = 'h60a6;
    'h2da : romdata_int = 'h278; // Line descriptor for 1_3
    'h2db : romdata_int = 'h4ccb;
    'h2dc : romdata_int = 'hb49;
    'h2dd : romdata_int = 'hef3;
    'h2de : romdata_int = 'h278; // Line descriptor for 1_3
    'h2df : romdata_int = 'h70b8;
    'h2e0 : romdata_int = 'h4a2c;
    'h2e1 : romdata_int = 'h4cee;
    'h2e2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2e3 : romdata_int = 'h2b8;
    'h2e4 : romdata_int = 'h4a5;
    'h2e5 : romdata_int = 'h341c;
    'h2e6 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h2e7 : romdata_int = 'h137;
    'h2e8 : romdata_int = 'h2687;
    'h2e9 : romdata_int = 'h5ab4;
    'h2ea : romdata_int = 'h278; // Line descriptor for 1_3
    'h2eb : romdata_int = 'h890;
    'h2ec : romdata_int = 'h1c78;
    'h2ed : romdata_int = 'h36ef;
    'h2ee : romdata_int = 'h278; // Line descriptor for 1_3
    'h2ef : romdata_int = 'h302;
    'h2f0 : romdata_int = 'h6665;
    'h2f1 : romdata_int = 'h72e1;
    'h2f2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2f3 : romdata_int = 'h3032;
    'h2f4 : romdata_int = 'h3e0d;
    'h2f5 : romdata_int = 'h4c4f;
    'h2f6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2f7 : romdata_int = 'h16ee;
    'h2f8 : romdata_int = 'h1a2c;
    'h2f9 : romdata_int = 'h1a9a;
    'h2fa : romdata_int = 'h4278; // Line descriptor for 1_3
    'h2fb : romdata_int = 'h251e;
    'h2fc : romdata_int = 'h473e;
    'h2fd : romdata_int = 'h6f0b;
    'h2fe : romdata_int = 'h278; // Line descriptor for 1_3
    'h2ff : romdata_int = 'hc9f;
    'h300 : romdata_int = 'h22c8;
    'h301 : romdata_int = 'h6325;
    'h302 : romdata_int = 'h278; // Line descriptor for 1_3
    'h303 : romdata_int = 'h263d;
    'h304 : romdata_int = 'h12c0;
    'h305 : romdata_int = 'h1218;
    'h306 : romdata_int = 'h278; // Line descriptor for 1_3
    'h307 : romdata_int = 'h1835;
    'h308 : romdata_int = 'h1882;
    'h309 : romdata_int = 'h26d9;
    'h30a : romdata_int = 'h278; // Line descriptor for 1_3
    'h30b : romdata_int = 'h62df;
    'h30c : romdata_int = 'h2759;
    'h30d : romdata_int = 'h263a;
    'h30e : romdata_int = 'h4278; // Line descriptor for 1_3
    'h30f : romdata_int = 'h467;
    'h310 : romdata_int = 'h6a7;
    'h311 : romdata_int = 'h12eb;
    'h312 : romdata_int = 'h278; // Line descriptor for 1_3
    'h313 : romdata_int = 'h5364;
    'h314 : romdata_int = 'h1ca6;
    'h315 : romdata_int = 'h395f;
    'h316 : romdata_int = 'h278; // Line descriptor for 1_3
    'h317 : romdata_int = 'he1a;
    'h318 : romdata_int = 'h12fd;
    'h319 : romdata_int = 'h5352;
    'h31a : romdata_int = 'h278; // Line descriptor for 1_3
    'h31b : romdata_int = 'h8;
    'h31c : romdata_int = 'h1ca8;
    'h31d : romdata_int = 'h4854;
    'h31e : romdata_int = 'h278; // Line descriptor for 1_3
    'h31f : romdata_int = 'h27f;
    'h320 : romdata_int = 'h3419;
    'h321 : romdata_int = 'h3cbd;
    'h322 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h323 : romdata_int = 'h147f;
    'h324 : romdata_int = 'h210b;
    'h325 : romdata_int = 'h3352;
    'h326 : romdata_int = 'h278; // Line descriptor for 1_3
    'h327 : romdata_int = 'hb27;
    'h328 : romdata_int = 'h1033;
    'h329 : romdata_int = 'h3e79;
    'h32a : romdata_int = 'h278; // Line descriptor for 1_3
    'h32b : romdata_int = 'h1b31;
    'h32c : romdata_int = 'hc70;
    'h32d : romdata_int = 'h8b6;
    'h32e : romdata_int = 'h278; // Line descriptor for 1_3
    'h32f : romdata_int = 'h4f4e;
    'h330 : romdata_int = 'h5e05;
    'h331 : romdata_int = 'h1a0a;
    'h332 : romdata_int = 'h278; // Line descriptor for 1_3
    'h333 : romdata_int = 'hc75;
    'h334 : romdata_int = 'h1208;
    'h335 : romdata_int = 'h550b;
    'h336 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h337 : romdata_int = 'h1050;
    'h338 : romdata_int = 'h1ac4;
    'h339 : romdata_int = 'h424f;
    'h33a : romdata_int = 'h278; // Line descriptor for 1_3
    'h33b : romdata_int = 'h67c;
    'h33c : romdata_int = 'h6a4;
    'h33d : romdata_int = 'hd38;
    'h33e : romdata_int = 'h278; // Line descriptor for 1_3
    'h33f : romdata_int = 'h3955;
    'h340 : romdata_int = 'h4134;
    'h341 : romdata_int = 'h5a38;
    'h342 : romdata_int = 'h278; // Line descriptor for 1_3
    'h343 : romdata_int = 'hc82;
    'h344 : romdata_int = 'h553d;
    'h345 : romdata_int = 'h6ef4;
    'h346 : romdata_int = 'h278; // Line descriptor for 1_3
    'h347 : romdata_int = 'h122;
    'h348 : romdata_int = 'h2126;
    'h349 : romdata_int = 'h50b3;
    'h34a : romdata_int = 'h4278; // Line descriptor for 1_3
    'h34b : romdata_int = 'h29b;
    'h34c : romdata_int = 'h105f;
    'h34d : romdata_int = 'h7015;
    'h34e : romdata_int = 'h278; // Line descriptor for 1_3
    'h34f : romdata_int = 'h125d;
    'h350 : romdata_int = 'h40d;
    'h351 : romdata_int = 'h27c;
    'h352 : romdata_int = 'h278; // Line descriptor for 1_3
    'h353 : romdata_int = 'h1873;
    'h354 : romdata_int = 'h2698;
    'h355 : romdata_int = 'h6944;
    'h356 : romdata_int = 'h278; // Line descriptor for 1_3
    'h357 : romdata_int = 'h127b;
    'h358 : romdata_int = 'h575c;
    'h359 : romdata_int = 'h1867;
    'h35a : romdata_int = 'h278; // Line descriptor for 1_3
    'h35b : romdata_int = 'h294c;
    'h35c : romdata_int = 'h5f25;
    'h35d : romdata_int = 'h74d9;
    'h35e : romdata_int = 'h4278; // Line descriptor for 1_3
    'h35f : romdata_int = 'h6a6;
    'h360 : romdata_int = 'h1ac9;
    'h361 : romdata_int = 'h2360;
    'h362 : romdata_int = 'h278; // Line descriptor for 1_3
    'h363 : romdata_int = 'heee;
    'h364 : romdata_int = 'h1e6b;
    'h365 : romdata_int = 'h6245;
    'h366 : romdata_int = 'h278; // Line descriptor for 1_3
    'h367 : romdata_int = 'h1d4b;
    'h368 : romdata_int = 'h2262;
    'h369 : romdata_int = 'h446b;
    'h36a : romdata_int = 'h278; // Line descriptor for 1_3
    'h36b : romdata_int = 'h8f2;
    'h36c : romdata_int = 'h271c;
    'h36d : romdata_int = 'h2721;
    'h36e : romdata_int = 'h278; // Line descriptor for 1_3
    'h36f : romdata_int = 'h2b44;
    'h370 : romdata_int = 'h3e81;
    'h371 : romdata_int = 'h214c;
    'h372 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h373 : romdata_int = 'h1b5b;
    'h374 : romdata_int = 'h5038;
    'h375 : romdata_int = 'h2a76;
    'h376 : romdata_int = 'h278; // Line descriptor for 1_3
    'h377 : romdata_int = 'h18c5;
    'h378 : romdata_int = 'h3d5b;
    'h379 : romdata_int = 'h6629;
    'h37a : romdata_int = 'h278; // Line descriptor for 1_3
    'h37b : romdata_int = 'h260;
    'h37c : romdata_int = 'ha48;
    'h37d : romdata_int = 'he0a;
    'h37e : romdata_int = 'h278; // Line descriptor for 1_3
    'h37f : romdata_int = 'h643;
    'h380 : romdata_int = 'h6b0;
    'h381 : romdata_int = 'h5506;
    'h382 : romdata_int = 'h278; // Line descriptor for 1_3
    'h383 : romdata_int = 'h238;
    'h384 : romdata_int = 'he32;
    'h385 : romdata_int = 'h10a2;
    'h386 : romdata_int = 'h6278; // Line descriptor for 1_3
    'h387 : romdata_int = 'h528;
    'h388 : romdata_int = 'h1cf5;
    'h389 : romdata_int = 'h492f;
    'h38a : romdata_int = 'h36c; // Line descriptor for 2_5
    'h38b : romdata_int = 'h2e;
    'h38c : romdata_int = 'hb0;
    'h38d : romdata_int = 'h4107;
    'h38e : romdata_int = 'h8f1c;
    'h38f : romdata_int = 'h36c; // Line descriptor for 2_5
    'h390 : romdata_int = 'h22f3;
    'h391 : romdata_int = 'h2680;
    'h392 : romdata_int = 'h2ead;
    'h393 : romdata_int = 'h5a42;
    'h394 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h395 : romdata_int = 'hd38;
    'h396 : romdata_int = 'h1763;
    'h397 : romdata_int = 'h38d6;
    'h398 : romdata_int = 'h5089;
    'h399 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h39a : romdata_int = 'h27f;
    'h39b : romdata_int = 'h1937;
    'h39c : romdata_int = 'h2ed5;
    'h39d : romdata_int = 'h632a;
    'h39e : romdata_int = 'h36c; // Line descriptor for 2_5
    'h39f : romdata_int = 'habd;
    'h3a0 : romdata_int = 'h1b4c;
    'h3a1 : romdata_int = 'h2107;
    'h3a2 : romdata_int = 'h8e89;
    'h3a3 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3a4 : romdata_int = 'h8c9;
    'h3a5 : romdata_int = 'ha67;
    'h3a6 : romdata_int = 'h1c14;
    'h3a7 : romdata_int = 'h853a;
    'h3a8 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3a9 : romdata_int = 'h14e5;
    'h3aa : romdata_int = 'h2236;
    'h3ab : romdata_int = 'h22f9;
    'h3ac : romdata_int = 'h5896;
    'h3ad : romdata_int = 'h436c; // Line descriptor for 2_5
    'h3ae : romdata_int = 'h1338;
    'h3af : romdata_int = 'h30a0;
    'h3b0 : romdata_int = 'h403d;
    'h3b1 : romdata_int = 'h7b3d;
    'h3b2 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3b3 : romdata_int = 'h10df;
    'h3b4 : romdata_int = 'h1887;
    'h3b5 : romdata_int = 'h28b1;
    'h3b6 : romdata_int = 'h5c58;
    'h3b7 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3b8 : romdata_int = 'h461;
    'h3b9 : romdata_int = 'h1408;
    'h3ba : romdata_int = 'h26db;
    'h3bb : romdata_int = 'h5718;
    'h3bc : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3bd : romdata_int = 'h1690;
    'h3be : romdata_int = 'h24e2;
    'h3bf : romdata_int = 'h2ae6;
    'h3c0 : romdata_int = 'h8663;
    'h3c1 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h3c2 : romdata_int = 'h183e;
    'h3c3 : romdata_int = 'h1ea6;
    'h3c4 : romdata_int = 'h226c;
    'h3c5 : romdata_int = 'h54a0;
    'h3c6 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3c7 : romdata_int = 'h86;
    'h3c8 : romdata_int = 'h4e0;
    'h3c9 : romdata_int = 'h2a26;
    'h3ca : romdata_int = 'h5ccb;
    'h3cb : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3cc : romdata_int = 'hf48;
    'h3cd : romdata_int = 'h89;
    'h3ce : romdata_int = 'h78cd;
    'h3cf : romdata_int = 'h1135;
    'h3d0 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3d1 : romdata_int = 'h1ced;
    'h3d2 : romdata_int = 'h3735;
    'h3d3 : romdata_int = 'h3521;
    'h3d4 : romdata_int = 'h5ed9;
    'h3d5 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h3d6 : romdata_int = 'h727a;
    'h3d7 : romdata_int = 'h1ccb;
    'h3d8 : romdata_int = 'h2d08;
    'h3d9 : romdata_int = 'h2f62;
    'h3da : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3db : romdata_int = 'h1ef5;
    'h3dc : romdata_int = 'h22ee;
    'h3dd : romdata_int = 'h7661;
    'h3de : romdata_int = 'h2aba;
    'h3df : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3e0 : romdata_int = 'h877;
    'h3e1 : romdata_int = 'h1144;
    'h3e2 : romdata_int = 'h2ee4;
    'h3e3 : romdata_int = 'h760b;
    'h3e4 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3e5 : romdata_int = 'hea1;
    'h3e6 : romdata_int = 'h12ce;
    'h3e7 : romdata_int = 'h2a70;
    'h3e8 : romdata_int = 'h7ec4;
    'h3e9 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h3ea : romdata_int = 'hd4f;
    'h3eb : romdata_int = 'h10d6;
    'h3ec : romdata_int = 'h1746;
    'h3ed : romdata_int = 'h887a;
    'h3ee : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3ef : romdata_int = 'h33b;
    'h3f0 : romdata_int = 'haa6;
    'h3f1 : romdata_int = 'h1b15;
    'h3f2 : romdata_int = 'h760e;
    'h3f3 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3f4 : romdata_int = 'hf2a;
    'h3f5 : romdata_int = 'h1d1f;
    'h3f6 : romdata_int = 'h2c0d;
    'h3f7 : romdata_int = 'h60ad;
    'h3f8 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3f9 : romdata_int = 'h46b;
    'h3fa : romdata_int = 'h18c3;
    'h3fb : romdata_int = 'h2034;
    'h3fc : romdata_int = 'h7046;
    'h3fd : romdata_int = 'h436c; // Line descriptor for 2_5
    'h3fe : romdata_int = 'h4;
    'h3ff : romdata_int = 'h12fe;
    'h400 : romdata_int = 'h145d;
    'h401 : romdata_int = 'h82b8;
    'h402 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h403 : romdata_int = 'h642;
    'h404 : romdata_int = 'h84a;
    'h405 : romdata_int = 'haf2;
    'h406 : romdata_int = 'h62fe;
    'h407 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h408 : romdata_int = 'h209e;
    'h409 : romdata_int = 'h267e;
    'h40a : romdata_int = 'h30b0;
    'h40b : romdata_int = 'h7062;
    'h40c : romdata_int = 'h36c; // Line descriptor for 2_5
    'h40d : romdata_int = 'h8d5;
    'h40e : romdata_int = 'h108d;
    'h40f : romdata_int = 'h2667;
    'h410 : romdata_int = 'h6b09;
    'h411 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h412 : romdata_int = 'h312;
    'h413 : romdata_int = 'h2039;
    'h414 : romdata_int = 'h2d1d;
    'h415 : romdata_int = 'h4eea;
    'h416 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h417 : romdata_int = 'hd4d;
    'h418 : romdata_int = 'h10a0;
    'h419 : romdata_int = 'h444b;
    'h41a : romdata_int = 'h6517;
    'h41b : romdata_int = 'h36c; // Line descriptor for 2_5
    'h41c : romdata_int = 'h299;
    'h41d : romdata_int = 'h92b;
    'h41e : romdata_int = 'h2e18;
    'h41f : romdata_int = 'h8149;
    'h420 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h421 : romdata_int = 'hcab;
    'h422 : romdata_int = 'h6703;
    'h423 : romdata_int = 'h6b0;
    'h424 : romdata_int = 'h2549;
    'h425 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h426 : romdata_int = 'h3762;
    'h427 : romdata_int = 'hc8f;
    'h428 : romdata_int = 'h6ab6;
    'h429 : romdata_int = 'h16b4;
    'h42a : romdata_int = 'h36c; // Line descriptor for 2_5
    'h42b : romdata_int = 'h1221;
    'h42c : romdata_int = 'h1e3f;
    'h42d : romdata_int = 'h2467;
    'h42e : romdata_int = 'h4c86;
    'h42f : romdata_int = 'h36c; // Line descriptor for 2_5
    'h430 : romdata_int = 'h3ed1;
    'h431 : romdata_int = 'h8b20;
    'h432 : romdata_int = 'h12fd;
    'h433 : romdata_int = 'h2291;
    'h434 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h435 : romdata_int = 'h9a;
    'h436 : romdata_int = 'h14c0;
    'h437 : romdata_int = 'h1f38;
    'h438 : romdata_int = 'h72f8;
    'h439 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h43a : romdata_int = 'hc70;
    'h43b : romdata_int = 'h1a64;
    'h43c : romdata_int = 'h2ae3;
    'h43d : romdata_int = 'h8706;
    'h43e : romdata_int = 'h36c; // Line descriptor for 2_5
    'h43f : romdata_int = 'h121c;
    'h440 : romdata_int = 'h1f4b;
    'h441 : romdata_int = 'h2257;
    'h442 : romdata_int = 'h6109;
    'h443 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h444 : romdata_int = 'h455;
    'h445 : romdata_int = 'h167e;
    'h446 : romdata_int = 'h430f;
    'h447 : romdata_int = 'h826b;
    'h448 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h449 : romdata_int = 'h109b;
    'h44a : romdata_int = 'h1b58;
    'h44b : romdata_int = 'h18ca;
    'h44c : romdata_int = 'h7c7b;
    'h44d : romdata_int = 'h436c; // Line descriptor for 2_5
    'h44e : romdata_int = 'h864;
    'h44f : romdata_int = 'h168f;
    'h450 : romdata_int = 'h1aad;
    'h451 : romdata_int = 'h4a4e;
    'h452 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h453 : romdata_int = 'he66;
    'h454 : romdata_int = 'h208b;
    'h455 : romdata_int = 'h6525;
    'h456 : romdata_int = 'h2c79;
    'h457 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h458 : romdata_int = 'h936;
    'h459 : romdata_int = 'ha88;
    'h45a : romdata_int = 'h26b5;
    'h45b : romdata_int = 'h6505;
    'h45c : romdata_int = 'h36c; // Line descriptor for 2_5
    'h45d : romdata_int = 'h2469;
    'h45e : romdata_int = 'hae;
    'h45f : romdata_int = 'h1b06;
    'h460 : romdata_int = 'h7553;
    'h461 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h462 : romdata_int = 'h1670;
    'h463 : romdata_int = 'h24ff;
    'h464 : romdata_int = 'h3326;
    'h465 : romdata_int = 'h88ca;
    'h466 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h467 : romdata_int = 'hf16;
    'h468 : romdata_int = 'h1ea1;
    'h469 : romdata_int = 'h2166;
    'h46a : romdata_int = 'h8a28;
    'h46b : romdata_int = 'h36c; // Line descriptor for 2_5
    'h46c : romdata_int = 'h4e6;
    'h46d : romdata_int = 'h161f;
    'h46e : romdata_int = 'h1a17;
    'h46f : romdata_int = 'h4af0;
    'h470 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h471 : romdata_int = 'hd5;
    'h472 : romdata_int = 'h2f3e;
    'h473 : romdata_int = 'h4009;
    'h474 : romdata_int = 'h7493;
    'h475 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h476 : romdata_int = 'hc41;
    'h477 : romdata_int = 'h1d3d;
    'h478 : romdata_int = 'h2630;
    'h479 : romdata_int = 'h88c3;
    'h47a : romdata_int = 'h36c; // Line descriptor for 2_5
    'h47b : romdata_int = 'h10b;
    'h47c : romdata_int = 'h51e;
    'h47d : romdata_int = 'h2b59;
    'h47e : romdata_int = 'h5248;
    'h47f : romdata_int = 'h36c; // Line descriptor for 2_5
    'h480 : romdata_int = 'h643;
    'h481 : romdata_int = 'h173f;
    'h482 : romdata_int = 'h293b;
    'h483 : romdata_int = 'h4a7b;
    'h484 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h485 : romdata_int = 'h2e54;
    'h486 : romdata_int = 'h6a7;
    'h487 : romdata_int = 'h687b;
    'h488 : romdata_int = 'h27c;
    'h489 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h48a : romdata_int = 'h44bb;
    'h48b : romdata_int = 'h5813;
    'h48c : romdata_int = 'h1a2b;
    'h48d : romdata_int = 'h6c9;
    'h48e : romdata_int = 'h36c; // Line descriptor for 2_5
    'h48f : romdata_int = 'h1319;
    'h490 : romdata_int = 'h1958;
    'h491 : romdata_int = 'h36e6;
    'h492 : romdata_int = 'h8a2c;
    'h493 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h494 : romdata_int = 'h22f4;
    'h495 : romdata_int = 'h2441;
    'h496 : romdata_int = 'h2c81;
    'h497 : romdata_int = 'h7d47;
    'h498 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h499 : romdata_int = 'hc0e;
    'h49a : romdata_int = 'h122a;
    'h49b : romdata_int = 'h1a42;
    'h49c : romdata_int = 'h4cb6;
    'h49d : romdata_int = 'h436c; // Line descriptor for 2_5
    'h49e : romdata_int = 'h10d0;
    'h49f : romdata_int = 'h255e;
    'h4a0 : romdata_int = 'h26a8;
    'h4a1 : romdata_int = 'h7260;
    'h4a2 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4a3 : romdata_int = 'he4d;
    'h4a4 : romdata_int = 'h1030;
    'h4a5 : romdata_int = 'h3270;
    'h4a6 : romdata_int = 'h6874;
    'h4a7 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4a8 : romdata_int = 'h18db;
    'h4a9 : romdata_int = 'h2145;
    'h4aa : romdata_int = 'h2d4c;
    'h4ab : romdata_int = 'h80a1;
    'h4ac : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4ad : romdata_int = 'h48a;
    'h4ae : romdata_int = 'h4d5;
    'h4af : romdata_int = 'h1522;
    'h4b0 : romdata_int = 'h5f38;
    'h4b1 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h4b2 : romdata_int = 'h12c9;
    'h4b3 : romdata_int = 'h1845;
    'h4b4 : romdata_int = 'h46f7;
    'h4b5 : romdata_int = 'h664e;
    'h4b6 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4b7 : romdata_int = 'h1623;
    'h4b8 : romdata_int = 'hb22;
    'h4b9 : romdata_int = 'h520b;
    'h4ba : romdata_int = 'h42b8;
    'h4bb : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4bc : romdata_int = 'h5d67;
    'h4bd : romdata_int = 'h28d4;
    'h4be : romdata_int = 'h168c;
    'h4bf : romdata_int = 'h1d1d;
    'h4c0 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4c1 : romdata_int = 'h862;
    'h4c2 : romdata_int = 'hc25;
    'h4c3 : romdata_int = 'h2ec7;
    'h4c4 : romdata_int = 'h50ec;
    'h4c5 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h4c6 : romdata_int = 'h253f;
    'h4c7 : romdata_int = 'h266e;
    'h4c8 : romdata_int = 'h2d61;
    'h4c9 : romdata_int = 'h8537;
    'h4ca : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4cb : romdata_int = 'ha5c;
    'h4cc : romdata_int = 'h5ab5;
    'h4cd : romdata_int = 'h954;
    'h4ce : romdata_int = 'h2645;
    'h4cf : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4d0 : romdata_int = 'h668d;
    'h4d1 : romdata_int = 'h214d;
    'h4d2 : romdata_int = 'hb49;
    'h4d3 : romdata_int = 'h3b4f;
    'h4d4 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4d5 : romdata_int = 'h673;
    'h4d6 : romdata_int = 'h187b;
    'h4d7 : romdata_int = 'h2081;
    'h4d8 : romdata_int = 'h74c6;
    'h4d9 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h4da : romdata_int = 'h2b8;
    'h4db : romdata_int = 'h10be;
    'h4dc : romdata_int = 'h3c01;
    'h4dd : romdata_int = 'h4913;
    'h4de : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4df : romdata_int = 'h890;
    'h4e0 : romdata_int = 'h2151;
    'h4e1 : romdata_int = 'h4220;
    'h4e2 : romdata_int = 'h551d;
    'h4e3 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4e4 : romdata_int = 'hef3;
    'h4e5 : romdata_int = 'h2665;
    'h4e6 : romdata_int = 'h4750;
    'h4e7 : romdata_int = 'h62d2;
    'h4e8 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4e9 : romdata_int = 'h27b;
    'h4ea : romdata_int = 'h1006;
    'h4eb : romdata_int = 'h2749;
    'h4ec : romdata_int = 'h5431;
    'h4ed : romdata_int = 'h436c; // Line descriptor for 2_5
    'h4ee : romdata_int = 'h137;
    'h4ef : romdata_int = 'h16da;
    'h4f0 : romdata_int = 'h2e36;
    'h4f1 : romdata_int = 'h6c29;
    'h4f2 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4f3 : romdata_int = 'h4a5;
    'h4f4 : romdata_int = 'h24a4;
    'h4f5 : romdata_int = 'h2aed;
    'h4f6 : romdata_int = 'h6e6e;
    'h4f7 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4f8 : romdata_int = 'h29b;
    'h4f9 : romdata_int = 'h1031;
    'h4fa : romdata_int = 'h28f3;
    'h4fb : romdata_int = 'h56fa;
    'h4fc : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4fd : romdata_int = 'h185c;
    'h4fe : romdata_int = 'h18ee;
    'h4ff : romdata_int = 'h3e87;
    'h500 : romdata_int = 'h6a17;
    'h501 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h502 : romdata_int = 'h2449;
    'h503 : romdata_int = 'h3a61;
    'h504 : romdata_int = 'h3c42;
    'h505 : romdata_int = 'h60a7;
    'h506 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h507 : romdata_int = 'h6e5;
    'h508 : romdata_int = 'h1efc;
    'h509 : romdata_int = 'h30fc;
    'h50a : romdata_int = 'h4d54;
    'h50b : romdata_int = 'h36c; // Line descriptor for 2_5
    'h50c : romdata_int = 'h2a85;
    'h50d : romdata_int = 'h2d2c;
    'h50e : romdata_int = 'h8c33;
    'h50f : romdata_int = 'h3f61;
    'h510 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h511 : romdata_int = 'h143f;
    'h512 : romdata_int = 'h1a35;
    'h513 : romdata_int = 'h1c9a;
    'h514 : romdata_int = 'h8c2c;
    'h515 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h516 : romdata_int = 'h6a6;
    'h517 : romdata_int = 'h1906;
    'h518 : romdata_int = 'h255d;
    'h519 : romdata_int = 'h8e9c;
    'h51a : romdata_int = 'h36c; // Line descriptor for 2_5
    'h51b : romdata_int = 'h467;
    'h51c : romdata_int = 'he1a;
    'h51d : romdata_int = 'hf58;
    'h51e : romdata_int = 'h7a2f;
    'h51f : romdata_int = 'h36c; // Line descriptor for 2_5
    'h520 : romdata_int = 'h1418;
    'h521 : romdata_int = 'h271e;
    'h522 : romdata_int = 'h2c4f;
    'h523 : romdata_int = 'h7e0d;
    'h524 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h525 : romdata_int = 'h283d;
    'h526 : romdata_int = 'h28d9;
    'h527 : romdata_int = 'h2f2f;
    'h528 : romdata_int = 'h4e43;
    'h529 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h52a : romdata_int = 'h8;
    'h52b : romdata_int = 'hb27;
    'h52c : romdata_int = 'h14eb;
    'h52d : romdata_int = 'h86b9;
    'h52e : romdata_int = 'h36c; // Line descriptor for 2_5
    'h52f : romdata_int = 'h238;
    'h530 : romdata_int = 'h283a;
    'h531 : romdata_int = 'h2959;
    'h532 : romdata_int = 'h6889;
    'h533 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h534 : romdata_int = 'h14fd;
    'h535 : romdata_int = 'hc82;
    'h536 : romdata_int = 'h24c8;
    'h537 : romdata_int = 'h8332;
    'h538 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h539 : romdata_int = 'h7951;
    'h53a : romdata_int = 'h1440;
    'h53b : romdata_int = 'h1e97;
    'h53c : romdata_int = 'h1d31;
    'h53d : romdata_int = 'h436c; // Line descriptor for 2_5
    'h53e : romdata_int = 'h230b;
    'h53f : romdata_int = 'h28ba;
    'h540 : romdata_int = 'h395f;
    'h541 : romdata_int = 'h8448;
    'h542 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h543 : romdata_int = 'h8b6;
    'h544 : romdata_int = 'h1233;
    'h545 : romdata_int = 'h3470;
    'h546 : romdata_int = 'h487d;
    'h547 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h548 : romdata_int = 'hc75;
    'h549 : romdata_int = 'h1465;
    'h54a : romdata_int = 'h6e4d;
    'h54b : romdata_int = 'h2efc;
    'h54c : romdata_int = 'h36c; // Line descriptor for 2_5
    'h54d : romdata_int = 'h72c;
    'h54e : romdata_int = 'hd52;
    'h54f : romdata_int = 'h1ed5;
    'h550 : romdata_int = 'h6f06;
    'h551 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h552 : romdata_int = 'h3d47;
    'h553 : romdata_int = 'h4845;
    'h554 : romdata_int = 'h67c;
    'h555 : romdata_int = 'h1cc4;
    'h556 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h557 : romdata_int = 'hb34;
    'h558 : romdata_int = 'h1250;
    'h559 : romdata_int = 'h32ee;
    'h55a : romdata_int = 'h6cf3;
    'h55b : romdata_int = 'h36c; // Line descriptor for 2_5
    'h55c : romdata_int = 'h122;
    'h55d : romdata_int = 'h2099;
    'h55e : romdata_int = 'h2cc6;
    'h55f : romdata_int = 'h8c12;
    'h560 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h561 : romdata_int = 'h302;
    'h562 : romdata_int = 'h1a73;
    'h563 : romdata_int = 'h2898;
    'h564 : romdata_int = 'h5b28;
    'h565 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h566 : romdata_int = 'h40d;
    'h567 : romdata_int = 'h147b;
    'h568 : romdata_int = 'h1c0a;
    'h569 : romdata_int = 'h791a;
    'h56a : romdata_int = 'h36c; // Line descriptor for 2_5
    'h56b : romdata_int = 'h2ef5;
    'h56c : romdata_int = 'h3544;
    'h56d : romdata_int = 'h3913;
    'h56e : romdata_int = 'h570b;
    'h56f : romdata_int = 'h36c; // Line descriptor for 2_5
    'h570 : romdata_int = 'h62d;
    'h571 : romdata_int = 'h2851;
    'h572 : romdata_int = 'h2ac2;
    'h573 : romdata_int = 'h7008;
    'h574 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h575 : romdata_int = 'heee;
    'h576 : romdata_int = 'h224a;
    'h577 : romdata_int = 'h46a6;
    'h578 : romdata_int = 'h7a68;
    'h579 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h57a : romdata_int = 'h1cc9;
    'h57b : romdata_int = 'h206b;
    'h57c : romdata_int = 'h2326;
    'h57d : romdata_int = 'h5144;
    'h57e : romdata_int = 'h36c; // Line descriptor for 2_5
    'h57f : romdata_int = 'h1eb1;
    'h580 : romdata_int = 'h8f2;
    'h581 : romdata_int = 'h3b3d;
    'h582 : romdata_int = 'h4e29;
    'h583 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h584 : romdata_int = 'h2b43;
    'h585 : romdata_int = 'h2356;
    'h586 : romdata_int = 'h5f4b;
    'h587 : romdata_int = 'h1ea8;
    'h588 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h589 : romdata_int = 'hb01;
    'h58a : romdata_int = 'h1d5b;
    'h58b : romdata_int = 'h291c;
    'h58c : romdata_int = 'h5878;
    'h58d : romdata_int = 'h436c; // Line descriptor for 2_5
    'h58e : romdata_int = 'h1ac5;
    'h58f : romdata_int = 'h2a1b;
    'h590 : romdata_int = 'h2ae4;
    'h591 : romdata_int = 'h6c39;
    'h592 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h593 : romdata_int = 'h2d34;
    'h594 : romdata_int = 'h279;
    'h595 : romdata_int = 'he0a;
    'h596 : romdata_int = 'h7d08;
    'h597 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h598 : romdata_int = 'h728;
    'h599 : romdata_int = 'h2cf2;
    'h59a : romdata_int = 'h4525;
    'h59b : romdata_int = 'h80d9;
    'h59c : romdata_int = 'h36c; // Line descriptor for 2_5
    'h59d : romdata_int = 'h2b9;
    'h59e : romdata_int = 'ha48;
    'h59f : romdata_int = 'h12a2;
    'h5a0 : romdata_int = 'h7e52;
    'h5a1 : romdata_int = 'h636c; // Line descriptor for 2_5
    'h5a2 : romdata_int = 'h528;
    'h5a3 : romdata_int = 'he32;
    'h5a4 : romdata_int = 'h1efe;
    'h5a5 : romdata_int = 'h5201;
    'h5a6 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5a7 : romdata_int = 'h352c;
    'h5a8 : romdata_int = 'h3703;
    'h5a9 : romdata_int = 'h3c43;
    'h5aa : romdata_int = 'h4800;
    'h5ab : romdata_int = 'h94b5;
    'h5ac : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5ad : romdata_int = 'h1432;
    'h5ae : romdata_int = 'h143d;
    'h5af : romdata_int = 'h291e;
    'h5b0 : romdata_int = 'h4a00;
    'h5b1 : romdata_int = 'h529a;
    'h5b2 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5b3 : romdata_int = 'h81f;
    'h5b4 : romdata_int = 'h200e;
    'h5b5 : romdata_int = 'h373e;
    'h5b6 : romdata_int = 'h4c00;
    'h5b7 : romdata_int = 'h668a;
    'h5b8 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5b9 : romdata_int = 'h506;
    'h5ba : romdata_int = 'hc45;
    'h5bb : romdata_int = 'h210b;
    'h5bc : romdata_int = 'h4e00;
    'h5bd : romdata_int = 'h8960;
    'h5be : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5bf : romdata_int = 'h133d;
    'h5c0 : romdata_int = 'h30ef;
    'h5c1 : romdata_int = 'h4224;
    'h5c2 : romdata_int = 'h5000;
    'h5c3 : romdata_int = 'ha516;
    'h5c4 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5c5 : romdata_int = 'h698;
    'h5c6 : romdata_int = 'h1afe;
    'h5c7 : romdata_int = 'h3088;
    'h5c8 : romdata_int = 'h3cd1;
    'h5c9 : romdata_int = 'h5200;
    'h5ca : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5cb : romdata_int = 'h1d1e;
    'h5cc : romdata_int = 'h2a67;
    'h5cd : romdata_int = 'h40ec;
    'h5ce : romdata_int = 'h5400;
    'h5cf : romdata_int = 'h9952;
    'h5d0 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5d1 : romdata_int = 'h87e;
    'h5d2 : romdata_int = 'h382c;
    'h5d3 : romdata_int = 'h4509;
    'h5d4 : romdata_int = 'h5600;
    'h5d5 : romdata_int = 'hb2d6;
    'h5d6 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5d7 : romdata_int = 'h214c;
    'h5d8 : romdata_int = 'h240f;
    'h5d9 : romdata_int = 'h3d29;
    'h5da : romdata_int = 'h5800;
    'h5db : romdata_int = 'hae31;
    'h5dc : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5dd : romdata_int = 'h2b55;
    'h5de : romdata_int = 'h3155;
    'h5df : romdata_int = 'h5a00;
    'h5e0 : romdata_int = 'h7528;
    'h5e1 : romdata_int = 'h9f61;
    'h5e2 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5e3 : romdata_int = 'h21c;
    'h5e4 : romdata_int = 'h88c;
    'h5e5 : romdata_int = 'hab0;
    'h5e6 : romdata_int = 'h4a01;
    'h5e7 : romdata_int = 'h5c00;
    'h5e8 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5e9 : romdata_int = 'h1115;
    'h5ea : romdata_int = 'h26c8;
    'h5eb : romdata_int = 'h2885;
    'h5ec : romdata_int = 'h40aa;
    'h5ed : romdata_int = 'h5e00;
    'h5ee : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5ef : romdata_int = 'h1f4d;
    'h5f0 : romdata_int = 'h344f;
    'h5f1 : romdata_int = 'h42b5;
    'h5f2 : romdata_int = 'h6000;
    'h5f3 : romdata_int = 'h9cc5;
    'h5f4 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5f5 : romdata_int = 'h1064;
    'h5f6 : romdata_int = 'h2091;
    'h5f7 : romdata_int = 'h5d3b;
    'h5f8 : romdata_int = 'h6200;
    'h5f9 : romdata_int = 'h84e7;
    'h5fa : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5fb : romdata_int = 'h1c;
    'h5fc : romdata_int = 'h24e2;
    'h5fd : romdata_int = 'h6400;
    'h5fe : romdata_int = 'h7e64;
    'h5ff : romdata_int = 'h8683;
    'h600 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h601 : romdata_int = 'h1aa6;
    'h602 : romdata_int = 'h2f4f;
    'h603 : romdata_int = 'h3cb8;
    'h604 : romdata_int = 'h6600;
    'h605 : romdata_int = 'h7f2b;
    'h606 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h607 : romdata_int = 'hc87;
    'h608 : romdata_int = 'h16ef;
    'h609 : romdata_int = 'h6800;
    'h60a : romdata_int = 'h767c;
    'h60b : romdata_int = 'h9255;
    'h60c : romdata_int = 'h45a; // Line descriptor for 1_2
    'h60d : romdata_int = 'h10ad;
    'h60e : romdata_int = 'h3636;
    'h60f : romdata_int = 'h6279;
    'h610 : romdata_int = 'h6a00;
    'h611 : romdata_int = 'h712e;
    'h612 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h613 : romdata_int = 'h1c6e;
    'h614 : romdata_int = 'h2e33;
    'h615 : romdata_int = 'h3311;
    'h616 : romdata_int = 'h6c00;
    'h617 : romdata_int = 'ha2a1;
    'h618 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h619 : romdata_int = 'h4c0;
    'h61a : romdata_int = 'h1e8b;
    'h61b : romdata_int = 'h38a0;
    'h61c : romdata_int = 'h4c72;
    'h61d : romdata_int = 'h6e00;
    'h61e : romdata_int = 'h45a; // Line descriptor for 1_2
    'h61f : romdata_int = 'h1632;
    'h620 : romdata_int = 'h2622;
    'h621 : romdata_int = 'h3f25;
    'h622 : romdata_int = 'h7000;
    'h623 : romdata_int = 'h945e;
    'h624 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h625 : romdata_int = 'h132;
    'h626 : romdata_int = 'h1017;
    'h627 : romdata_int = 'h16bc;
    'h628 : romdata_int = 'h7200;
    'h629 : romdata_int = 'h8718;
    'h62a : romdata_int = 'h45a; // Line descriptor for 1_2
    'h62b : romdata_int = 'h2659;
    'h62c : romdata_int = 'h3f32;
    'h62d : romdata_int = 'h7400;
    'h62e : romdata_int = 'h8f22;
    'h62f : romdata_int = 'haa37;
    'h630 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h631 : romdata_int = 'h6cf;
    'h632 : romdata_int = 'h122c;
    'h633 : romdata_int = 'h26aa;
    'h634 : romdata_int = 'h5ab8;
    'h635 : romdata_int = 'h7600;
    'h636 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h637 : romdata_int = 'h823;
    'h638 : romdata_int = 'h2249;
    'h639 : romdata_int = 'h46cc;
    'h63a : romdata_int = 'h6861;
    'h63b : romdata_int = 'h7800;
    'h63c : romdata_int = 'h45a; // Line descriptor for 1_2
    'h63d : romdata_int = 'h2603;
    'h63e : romdata_int = 'h3121;
    'h63f : romdata_int = 'h36e4;
    'h640 : romdata_int = 'h7a00;
    'h641 : romdata_int = 'h9c4c;
    'h642 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h643 : romdata_int = 'h521;
    'h644 : romdata_int = 'h3a75;
    'h645 : romdata_int = 'h6855;
    'h646 : romdata_int = 'h7c00;
    'h647 : romdata_int = 'ha6f3;
    'h648 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h649 : romdata_int = 'he82;
    'h64a : romdata_int = 'h1aa8;
    'h64b : romdata_int = 'h4445;
    'h64c : romdata_int = 'h7e00;
    'h64d : romdata_int = 'h8413;
    'h64e : romdata_int = 'h45a; // Line descriptor for 1_2
    'h64f : romdata_int = 'h2511;
    'h650 : romdata_int = 'h334c;
    'h651 : romdata_int = 'h400a;
    'h652 : romdata_int = 'h5a7b;
    'h653 : romdata_int = 'h8000;
    'h654 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h655 : romdata_int = 'haee;
    'h656 : romdata_int = 'hcee;
    'h657 : romdata_int = 'h1c4a;
    'h658 : romdata_int = 'h468d;
    'h659 : romdata_int = 'h8200;
    'h65a : romdata_int = 'h45a; // Line descriptor for 1_2
    'h65b : romdata_int = 'h287e;
    'h65c : romdata_int = 'h2c3d;
    'h65d : romdata_int = 'h5e9b;
    'h65e : romdata_int = 'h8400;
    'h65f : romdata_int = 'hac1e;
    'h660 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h661 : romdata_int = 'h680;
    'h662 : romdata_int = 'h946;
    'h663 : romdata_int = 'h5cb9;
    'h664 : romdata_int = 'h8600;
    'h665 : romdata_int = 'ha0e9;
    'h666 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h667 : romdata_int = 'hcca;
    'h668 : romdata_int = 'h2349;
    'h669 : romdata_int = 'h32bd;
    'h66a : romdata_int = 'h80d5;
    'h66b : romdata_int = 'h8800;
    'h66c : romdata_int = 'h45a; // Line descriptor for 1_2
    'h66d : romdata_int = 'h1e6f;
    'h66e : romdata_int = 'h2057;
    'h66f : romdata_int = 'h4725;
    'h670 : romdata_int = 'h502e;
    'h671 : romdata_int = 'h8a00;
    'h672 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h673 : romdata_int = 'h162f;
    'h674 : romdata_int = 'h1920;
    'h675 : romdata_int = 'h8c00;
    'h676 : romdata_int = 'h9aab;
    'h677 : romdata_int = 'hb144;
    'h678 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h679 : romdata_int = 'h1ce5;
    'h67a : romdata_int = 'h2c98;
    'h67b : romdata_int = 'h38ad;
    'h67c : romdata_int = 'h4915;
    'h67d : romdata_int = 'h8e00;
    'h67e : romdata_int = 'h45a; // Line descriptor for 1_2
    'h67f : romdata_int = 'ha23;
    'h680 : romdata_int = 'h2ae5;
    'h681 : romdata_int = 'h3315;
    'h682 : romdata_int = 'h6728;
    'h683 : romdata_int = 'h9000;
    'h684 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h685 : romdata_int = 'h890;
    'h686 : romdata_int = 'h151d;
    'h687 : romdata_int = 'h3e45;
    'h688 : romdata_int = 'h7ac4;
    'h689 : romdata_int = 'h9200;
    'h68a : romdata_int = 'h45a; // Line descriptor for 1_2
    'h68b : romdata_int = 'he67;
    'h68c : romdata_int = 'h14a4;
    'h68d : romdata_int = 'h4a2b;
    'h68e : romdata_int = 'h642a;
    'h68f : romdata_int = 'h9400;
    'h690 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h691 : romdata_int = 'h2865;
    'h692 : romdata_int = 'h354c;
    'h693 : romdata_int = 'h6165;
    'h694 : romdata_int = 'h9600;
    'h695 : romdata_int = 'h6e5f;
    'h696 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h697 : romdata_int = 'h1f51;
    'h698 : romdata_int = 'h2858;
    'h699 : romdata_int = 'h8c88;
    'h69a : romdata_int = 'h9670;
    'h69b : romdata_int = 'h9800;
    'h69c : romdata_int = 'h45a; // Line descriptor for 1_2
    'h69d : romdata_int = 'h235d;
    'h69e : romdata_int = 'h3f13;
    'h69f : romdata_int = 'h72a7;
    'h6a0 : romdata_int = 'h7443;
    'h6a1 : romdata_int = 'h9a00;
    'h6a2 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6a3 : romdata_int = 'h2137;
    'h6a4 : romdata_int = 'h28ee;
    'h6a5 : romdata_int = 'h36f5;
    'h6a6 : romdata_int = 'h9c00;
    'h6a7 : romdata_int = 'hac49;
    'h6a8 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6a9 : romdata_int = 'h1c3c;
    'h6aa : romdata_int = 'h2a32;
    'h6ab : romdata_int = 'h7673;
    'h6ac : romdata_int = 'h9e00;
    'h6ad : romdata_int = 'hb2df;
    'h6ae : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6af : romdata_int = 'h103c;
    'h6b0 : romdata_int = 'h2694;
    'h6b1 : romdata_int = 'h326b;
    'h6b2 : romdata_int = 'h4e08;
    'h6b3 : romdata_int = 'ha000;
    'h6b4 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6b5 : romdata_int = 'h233;
    'h6b6 : romdata_int = 'ha44;
    'h6b7 : romdata_int = 'h243a;
    'h6b8 : romdata_int = 'h2cb1;
    'h6b9 : romdata_int = 'ha200;
    'h6ba : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6bb : romdata_int = 'he41;
    'h6bc : romdata_int = 'h2b49;
    'h6bd : romdata_int = 'h4219;
    'h6be : romdata_int = 'h8e48;
    'h6bf : romdata_int = 'ha400;
    'h6c0 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6c1 : romdata_int = 'h5f;
    'h6c2 : romdata_int = 'h34a5;
    'h6c3 : romdata_int = 'h64ef;
    'h6c4 : romdata_int = 'h8354;
    'h6c5 : romdata_int = 'ha600;
    'h6c6 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6c7 : romdata_int = 'h67;
    'h6c8 : romdata_int = 'h14b3;
    'h6c9 : romdata_int = 'h1ccc;
    'h6ca : romdata_int = 'h46d3;
    'h6cb : romdata_int = 'ha800;
    'h6cc : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6cd : romdata_int = 'h71;
    'h6ce : romdata_int = 'haba;
    'h6cf : romdata_int = 'h3a13;
    'h6d0 : romdata_int = 'h4328;
    'h6d1 : romdata_int = 'haa00;
    'h6d2 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6d3 : romdata_int = 'h338;
    'h6d4 : romdata_int = 'h16f8;
    'h6d5 : romdata_int = 'h1874;
    'h6d6 : romdata_int = 'h7894;
    'h6d7 : romdata_int = 'hac00;
    'h6d8 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6d9 : romdata_int = 'h228;
    'h6da : romdata_int = 'h640;
    'h6db : romdata_int = 'h2af3;
    'h6dc : romdata_int = 'hae00;
    'h6dd : romdata_int = 'haae5;
    'h6de : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6df : romdata_int = 'haeb;
    'h6e0 : romdata_int = 'h235e;
    'h6e1 : romdata_int = 'h932b;
    'h6e2 : romdata_int = 'hae8d;
    'h6e3 : romdata_int = 'hb000;
    'h6e4 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6e5 : romdata_int = 'h14f6;
    'h6e6 : romdata_int = 'h2e91;
    'h6e7 : romdata_int = 'h5089;
    'h6e8 : romdata_int = 'h88c5;
    'h6e9 : romdata_int = 'hb200;
    'h6ea : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6eb : romdata_int = 'h0;
    'h6ec : romdata_int = 'h722;
    'h6ed : romdata_int = 'hc5c;
    'h6ee : romdata_int = 'h1106;
    'h6ef : romdata_int = 'ha632;
    'h6f0 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6f1 : romdata_int = 'h200;
    'h6f2 : romdata_int = 'h335b;
    'h6f3 : romdata_int = 'h3c05;
    'h6f4 : romdata_int = 'h6aa5;
    'h6f5 : romdata_int = 'hb006;
    'h6f6 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6f7 : romdata_int = 'h400;
    'h6f8 : romdata_int = 'hd58;
    'h6f9 : romdata_int = 'h38b0;
    'h6fa : romdata_int = 'h3c20;
    'h6fb : romdata_int = 'h540b;
    'h6fc : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6fd : romdata_int = 'h600;
    'h6fe : romdata_int = 'h6ab;
    'h6ff : romdata_int = 'h186a;
    'h700 : romdata_int = 'h3534;
    'h701 : romdata_int = 'h786a;
    'h702 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h703 : romdata_int = 'h800;
    'h704 : romdata_int = 'h93f;
    'h705 : romdata_int = 'h3a38;
    'h706 : romdata_int = 'h2ecf;
    'h707 : romdata_int = 'h4717;
    'h708 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h709 : romdata_int = 'ha00;
    'h70a : romdata_int = 'h2269;
    'h70b : romdata_int = 'h3a70;
    'h70c : romdata_int = 'h5859;
    'h70d : romdata_int = 'h6cae;
    'h70e : romdata_int = 'h45a; // Line descriptor for 1_2
    'h70f : romdata_int = 'hc00;
    'h710 : romdata_int = 'h1967;
    'h711 : romdata_int = 'h2b37;
    'h712 : romdata_int = 'h4c02;
    'h713 : romdata_int = 'h732c;
    'h714 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h715 : romdata_int = 'he00;
    'h716 : romdata_int = 'h1956;
    'h717 : romdata_int = 'h3edf;
    'h718 : romdata_int = 'h7a4e;
    'h719 : romdata_int = 'h8d27;
    'h71a : romdata_int = 'h45a; // Line descriptor for 1_2
    'h71b : romdata_int = 'h1000;
    'h71c : romdata_int = 'h181e;
    'h71d : romdata_int = 'h1844;
    'h71e : romdata_int = 'h4662;
    'h71f : romdata_int = 'h82c9;
    'h720 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h721 : romdata_int = 'h221;
    'h722 : romdata_int = 'h250;
    'h723 : romdata_int = 'h1200;
    'h724 : romdata_int = 'h3b44;
    'h725 : romdata_int = 'h4484;
    'h726 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h727 : romdata_int = 'h6b4;
    'h728 : romdata_int = 'h1400;
    'h729 : romdata_int = 'h2447;
    'h72a : romdata_int = 'h2f44;
    'h72b : romdata_int = 'h42e1;
    'h72c : romdata_int = 'h45a; // Line descriptor for 1_2
    'h72d : romdata_int = 'h1600;
    'h72e : romdata_int = 'h1ad5;
    'h72f : romdata_int = 'h2267;
    'h730 : romdata_int = 'h5f12;
    'h731 : romdata_int = 'h9122;
    'h732 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h733 : romdata_int = 'hefd;
    'h734 : romdata_int = 'h1800;
    'h735 : romdata_int = 'h1e34;
    'h736 : romdata_int = 'h315f;
    'h737 : romdata_int = 'ha24d;
    'h738 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h739 : romdata_int = 'h12f6;
    'h73a : romdata_int = 'h1a00;
    'h73b : romdata_int = 'h3d0f;
    'h73c : romdata_int = 'h44e8;
    'h73d : romdata_int = 'h621e;
    'h73e : romdata_int = 'h45a; // Line descriptor for 1_2
    'h73f : romdata_int = 'hcc3;
    'h740 : romdata_int = 'h1c00;
    'h741 : romdata_int = 'h3ef7;
    'h742 : romdata_int = 'h40ce;
    'h743 : romdata_int = 'h563a;
    'h744 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h745 : romdata_int = 'h1e00;
    'h746 : romdata_int = 'h2d59;
    'h747 : romdata_int = 'h347e;
    'h748 : romdata_int = 'h9e8a;
    'h749 : romdata_int = 'ha858;
    'h74a : romdata_int = 'h45a; // Line descriptor for 1_2
    'h74b : romdata_int = 'h308;
    'h74c : romdata_int = 'h1af5;
    'h74d : romdata_int = 'h2000;
    'h74e : romdata_int = 'h2810;
    'h74f : romdata_int = 'h4089;
    'h750 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h751 : romdata_int = 'h512;
    'h752 : romdata_int = 'h2200;
    'h753 : romdata_int = 'h22a4;
    'h754 : romdata_int = 'h311c;
    'h755 : romdata_int = 'h383e;
    'h756 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h757 : romdata_int = 'h2400;
    'h758 : romdata_int = 'h408;
    'h759 : romdata_int = 'h44ad;
    'h75a : romdata_int = 'h4f0b;
    'h75b : romdata_int = 'h6ae0;
    'h75c : romdata_int = 'h45a; // Line descriptor for 1_2
    'h75d : romdata_int = 'h24b8;
    'h75e : romdata_int = 'h2600;
    'h75f : romdata_int = 'h374a;
    'h760 : romdata_int = 'h464e;
    'h761 : romdata_int = 'h7cd8;
    'h762 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h763 : romdata_int = 'h2d1c;
    'h764 : romdata_int = 'h1331;
    'h765 : romdata_int = 'h12bb;
    'h766 : romdata_int = 'h2800;
    'h767 : romdata_int = 'h9682;
    'h768 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h769 : romdata_int = 'h2a00;
    'h76a : romdata_int = 'h2cd9;
    'h76b : romdata_int = 'h2f60;
    'h76c : romdata_int = 'h8a67;
    'h76d : romdata_int = 'h9a0e;
    'h76e : romdata_int = 'h45a; // Line descriptor for 1_2
    'h76f : romdata_int = 'h1ccb;
    'h770 : romdata_int = 'h2c00;
    'h771 : romdata_int = 'h34f2;
    'h772 : romdata_int = 'h3b21;
    'h773 : romdata_int = 'h6d11;
    'h774 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h775 : romdata_int = 'he7d;
    'h776 : romdata_int = 'h2e00;
    'h777 : romdata_int = 'h3100;
    'h778 : romdata_int = 'h38fc;
    'h779 : romdata_int = 'h48a1;
    'h77a : romdata_int = 'h45a; // Line descriptor for 1_2
    'h77b : romdata_int = 'h1a97;
    'h77c : romdata_int = 'h1f13;
    'h77d : romdata_int = 'h3000;
    'h77e : romdata_int = 'h52b0;
    'h77f : romdata_int = 'h5938;
    'h780 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h781 : romdata_int = 'h465;
    'h782 : romdata_int = 'h2cf3;
    'h783 : romdata_int = 'h3200;
    'h784 : romdata_int = 'h60c7;
    'h785 : romdata_int = 'ha40a;
    'h786 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h787 : romdata_int = 'h43f;
    'h788 : romdata_int = 'h1b4b;
    'h789 : romdata_int = 'h3400;
    'h78a : romdata_int = 'h8062;
    'h78b : romdata_int = 'ha164;
    'h78c : romdata_int = 'h45a; // Line descriptor for 1_2
    'h78d : romdata_int = 'h20f3;
    'h78e : romdata_int = 'h3600;
    'h78f : romdata_int = 'h44fd;
    'h790 : romdata_int = 'h907c;
    'h791 : romdata_int = 'h994d;
    'h792 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h793 : romdata_int = 'h9f;
    'h794 : romdata_int = 'h131f;
    'h795 : romdata_int = 'h3800;
    'h796 : romdata_int = 'h44a7;
    'h797 : romdata_int = 'h6f62;
    'h798 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h799 : romdata_int = 'he9d;
    'h79a : romdata_int = 'h3602;
    'h79b : romdata_int = 'h3a00;
    'h79c : romdata_int = 'h42d9;
    'h79d : romdata_int = 'h7c0f;
    'h79e : romdata_int = 'h45a; // Line descriptor for 1_2
    'h79f : romdata_int = 'h16bd;
    'h7a0 : romdata_int = 'h2406;
    'h7a1 : romdata_int = 'h38f2;
    'h7a2 : romdata_int = 'h3c00;
    'h7a3 : romdata_int = 'h8b49;
    'h7a4 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h7a5 : romdata_int = 'h12ed;
    'h7a6 : romdata_int = 'h14a2;
    'h7a7 : romdata_int = 'h3e00;
    'h7a8 : romdata_int = 'h3b4e;
    'h7a9 : romdata_int = 'h4242;
    'h7aa : romdata_int = 'h45a; // Line descriptor for 1_2
    'h7ab : romdata_int = 'h114c;
    'h7ac : romdata_int = 'h2e76;
    'h7ad : romdata_int = 'h3f50;
    'h7ae : romdata_int = 'h4000;
    'h7af : romdata_int = 'h4144;
    'h7b0 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h7b1 : romdata_int = 'h1703;
    'h7b2 : romdata_int = 'h3361;
    'h7b3 : romdata_int = 'h4200;
    'h7b4 : romdata_int = 'h54ec;
    'h7b5 : romdata_int = 'ha8f1;
    'h7b6 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h7b7 : romdata_int = 'hab1;
    'h7b8 : romdata_int = 'he07;
    'h7b9 : romdata_int = 'h1e99;
    'h7ba : romdata_int = 'h4400;
    'h7bb : romdata_int = 'h70dd;
    'h7bc : romdata_int = 'h645a; // Line descriptor for 1_2
    'h7bd : romdata_int = 'h12a;
    'h7be : romdata_int = 'h26d8;
    'h7bf : romdata_int = 'h4166;
    'h7c0 : romdata_int = 'h4600;
    'h7c1 : romdata_int = 'h56a1;
    'h7c2 : romdata_int = 'h848; // Line descriptor for 3_5
    'h7c3 : romdata_int = 'hed;
    'h7c4 : romdata_int = 'h1ec8;
    'h7c5 : romdata_int = 'h2d39;
    'h7c6 : romdata_int = 'h3086;
    'h7c7 : romdata_int = 'h4159;
    'h7c8 : romdata_int = 'h4272;
    'h7c9 : romdata_int = 'h4800;
    'h7ca : romdata_int = 'h50d1;
    'h7cb : romdata_int = 'hcacb;
    'h7cc : romdata_int = 'h4848; // Line descriptor for 3_5
    'h7cd : romdata_int = 'h9b;
    'h7ce : romdata_int = 'he8a;
    'h7cf : romdata_int = 'h121a;
    'h7d0 : romdata_int = 'h1706;
    'h7d1 : romdata_int = 'h3043;
    'h7d2 : romdata_int = 'h4286;
    'h7d3 : romdata_int = 'h4a00;
    'h7d4 : romdata_int = 'h584a;
    'h7d5 : romdata_int = 'hc35a;
    'h7d6 : romdata_int = 'h848; // Line descriptor for 3_5
    'h7d7 : romdata_int = 'h565;
    'h7d8 : romdata_int = 'hd01;
    'h7d9 : romdata_int = 'h10b2;
    'h7da : romdata_int = 'h1c34;
    'h7db : romdata_int = 'h429c;
    'h7dc : romdata_int = 'h4423;
    'h7dd : romdata_int = 'h4c00;
    'h7de : romdata_int = 'h805e;
    'h7df : romdata_int = 'hb953;
    'h7e0 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h7e1 : romdata_int = 'h1947;
    'h7e2 : romdata_int = 'h22ba;
    'h7e3 : romdata_int = 'h22d9;
    'h7e4 : romdata_int = 'h2c91;
    'h7e5 : romdata_int = 'h3503;
    'h7e6 : romdata_int = 'h36f3;
    'h7e7 : romdata_int = 'h4e00;
    'h7e8 : romdata_int = 'h7367;
    'h7e9 : romdata_int = 'hd0d3;
    'h7ea : romdata_int = 'h848; // Line descriptor for 3_5
    'h7eb : romdata_int = 'hf61;
    'h7ec : romdata_int = 'h167d;
    'h7ed : romdata_int = 'h1c8b;
    'h7ee : romdata_int = 'h2432;
    'h7ef : romdata_int = 'h2479;
    'h7f0 : romdata_int = 'h3222;
    'h7f1 : romdata_int = 'h5000;
    'h7f2 : romdata_int = 'h6e17;
    'h7f3 : romdata_int = 'hc166;
    'h7f4 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h7f5 : romdata_int = 'h2cd1;
    'h7f6 : romdata_int = 'h30d2;
    'h7f7 : romdata_int = 'h32a0;
    'h7f8 : romdata_int = 'h380b;
    'h7f9 : romdata_int = 'h3a35;
    'h7fa : romdata_int = 'h3e78;
    'h7fb : romdata_int = 'h5200;
    'h7fc : romdata_int = 'h60c9;
    'h7fd : romdata_int = 'hbc89;
    'h7fe : romdata_int = 'h848; // Line descriptor for 3_5
    'h7ff : romdata_int = 'hc55;
    'h800 : romdata_int = 'h14b4;
    'h801 : romdata_int = 'h1864;
    'h802 : romdata_int = 'h2360;
    'h803 : romdata_int = 'h28f5;
    'h804 : romdata_int = 'h331d;
    'h805 : romdata_int = 'h5400;
    'h806 : romdata_int = 'h64b8;
    'h807 : romdata_int = 'hc555;
    'h808 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h809 : romdata_int = 'h143e;
    'h80a : romdata_int = 'h24e4;
    'h80b : romdata_int = 'h32b8;
    'h80c : romdata_int = 'h372a;
    'h80d : romdata_int = 'h3c56;
    'h80e : romdata_int = 'h3e2c;
    'h80f : romdata_int = 'h5600;
    'h810 : romdata_int = 'h5b03;
    'h811 : romdata_int = 'hc31f;
    'h812 : romdata_int = 'h848; // Line descriptor for 3_5
    'h813 : romdata_int = 'h762;
    'h814 : romdata_int = 'h1062;
    'h815 : romdata_int = 'h1058;
    'h816 : romdata_int = 'h1079;
    'h817 : romdata_int = 'h2c38;
    'h818 : romdata_int = 'h46f6;
    'h819 : romdata_int = 'h4c82;
    'h81a : romdata_int = 'h5800;
    'h81b : romdata_int = 'h9f65;
    'h81c : romdata_int = 'h4848; // Line descriptor for 3_5
    'h81d : romdata_int = 'h4e;
    'h81e : romdata_int = 'he75;
    'h81f : romdata_int = 'h169d;
    'h820 : romdata_int = 'h2c42;
    'h821 : romdata_int = 'h3d49;
    'h822 : romdata_int = 'h3ea9;
    'h823 : romdata_int = 'h5a00;
    'h824 : romdata_int = 'h8640;
    'h825 : romdata_int = 'h9b56;
    'h826 : romdata_int = 'h848; // Line descriptor for 3_5
    'h827 : romdata_int = 'h23a;
    'h828 : romdata_int = 'h1a3d;
    'h829 : romdata_int = 'h2251;
    'h82a : romdata_int = 'h2ebb;
    'h82b : romdata_int = 'h30ea;
    'h82c : romdata_int = 'h3c83;
    'h82d : romdata_int = 'h5c00;
    'h82e : romdata_int = 'h670b;
    'h82f : romdata_int = 'hce0d;
    'h830 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h831 : romdata_int = 'h86a;
    'h832 : romdata_int = 'h132c;
    'h833 : romdata_int = 'h165c;
    'h834 : romdata_int = 'h1688;
    'h835 : romdata_int = 'h1f50;
    'h836 : romdata_int = 'h20f3;
    'h837 : romdata_int = 'h5e00;
    'h838 : romdata_int = 'h703d;
    'h839 : romdata_int = 'ha520;
    'h83a : romdata_int = 'h848; // Line descriptor for 3_5
    'h83b : romdata_int = 'ha4a;
    'h83c : romdata_int = 'h16ca;
    'h83d : romdata_int = 'h1aa2;
    'h83e : romdata_int = 'h3318;
    'h83f : romdata_int = 'h435a;
    'h840 : romdata_int = 'h4667;
    'h841 : romdata_int = 'h5300;
    'h842 : romdata_int = 'h6000;
    'h843 : romdata_int = 'hbc72;
    'h844 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h845 : romdata_int = 'h65f;
    'h846 : romdata_int = 'h6dd;
    'h847 : romdata_int = 'he33;
    'h848 : romdata_int = 'h1f3f;
    'h849 : romdata_int = 'h3e28;
    'h84a : romdata_int = 'h44a3;
    'h84b : romdata_int = 'h4903;
    'h84c : romdata_int = 'h6200;
    'h84d : romdata_int = 'ha20e;
    'h84e : romdata_int = 'h848; // Line descriptor for 3_5
    'h84f : romdata_int = 'he41;
    'h850 : romdata_int = 'h1b1d;
    'h851 : romdata_int = 'h1e6f;
    'h852 : romdata_int = 'h234c;
    'h853 : romdata_int = 'h393e;
    'h854 : romdata_int = 'h3b60;
    'h855 : romdata_int = 'h6400;
    'h856 : romdata_int = 'h8a1c;
    'h857 : romdata_int = 'hb260;
    'h858 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h859 : romdata_int = 'h8c9;
    'h85a : romdata_int = 'h1e69;
    'h85b : romdata_int = 'h2f32;
    'h85c : romdata_int = 'h36e2;
    'h85d : romdata_int = 'h3e8f;
    'h85e : romdata_int = 'h4075;
    'h85f : romdata_int = 'h6600;
    'h860 : romdata_int = 'h78df;
    'h861 : romdata_int = 'ha0a7;
    'h862 : romdata_int = 'h848; // Line descriptor for 3_5
    'h863 : romdata_int = 'h1341;
    'h864 : romdata_int = 'h1af6;
    'h865 : romdata_int = 'h1e47;
    'h866 : romdata_int = 'h2700;
    'h867 : romdata_int = 'h3706;
    'h868 : romdata_int = 'h3a46;
    'h869 : romdata_int = 'h5356;
    'h86a : romdata_int = 'h6800;
    'h86b : romdata_int = 'hcc33;
    'h86c : romdata_int = 'h4848; // Line descriptor for 3_5
    'h86d : romdata_int = 'h41e;
    'h86e : romdata_int = 'hb60;
    'h86f : romdata_int = 'h2e05;
    'h870 : romdata_int = 'h34cc;
    'h871 : romdata_int = 'h3b3f;
    'h872 : romdata_int = 'h4658;
    'h873 : romdata_int = 'h6a00;
    'h874 : romdata_int = 'h792c;
    'h875 : romdata_int = 'hb456;
    'h876 : romdata_int = 'h848; // Line descriptor for 3_5
    'h877 : romdata_int = 'h2e1;
    'h878 : romdata_int = 'h8f2;
    'h879 : romdata_int = 'h1c28;
    'h87a : romdata_int = 'h1c81;
    'h87b : romdata_int = 'h2854;
    'h87c : romdata_int = 'h2f50;
    'h87d : romdata_int = 'h6c00;
    'h87e : romdata_int = 'h753c;
    'h87f : romdata_int = 'hc6ac;
    'h880 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h881 : romdata_int = 'h4bc;
    'h882 : romdata_int = 'ha4e;
    'h883 : romdata_int = 'hf64;
    'h884 : romdata_int = 'h1268;
    'h885 : romdata_int = 'h3629;
    'h886 : romdata_int = 'h3e33;
    'h887 : romdata_int = 'h6e00;
    'h888 : romdata_int = 'h76c4;
    'h889 : romdata_int = 'hb6c1;
    'h88a : romdata_int = 'h848; // Line descriptor for 3_5
    'h88b : romdata_int = 'h479;
    'h88c : romdata_int = 'h1522;
    'h88d : romdata_int = 'h1733;
    'h88e : romdata_int = 'h267a;
    'h88f : romdata_int = 'h2ea6;
    'h890 : romdata_int = 'h4130;
    'h891 : romdata_int = 'h7000;
    'h892 : romdata_int = 'h7e70;
    'h893 : romdata_int = 'hb8b7;
    'h894 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h895 : romdata_int = 'h50b;
    'h896 : romdata_int = 'h6e6;
    'h897 : romdata_int = 'h950;
    'h898 : romdata_int = 'hc4b;
    'h899 : romdata_int = 'h1eb5;
    'h89a : romdata_int = 'h24e3;
    'h89b : romdata_int = 'h7200;
    'h89c : romdata_int = 'h7c08;
    'h89d : romdata_int = 'h9647;
    'h89e : romdata_int = 'h848; // Line descriptor for 3_5
    'h89f : romdata_int = 'h72e;
    'h8a0 : romdata_int = 'h223a;
    'h8a1 : romdata_int = 'h2ae6;
    'h8a2 : romdata_int = 'h348d;
    'h8a3 : romdata_int = 'h34d3;
    'h8a4 : romdata_int = 'h3b08;
    'h8a5 : romdata_int = 'h620a;
    'h8a6 : romdata_int = 'h7400;
    'h8a7 : romdata_int = 'hccec;
    'h8a8 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h8a9 : romdata_int = 'h2ec;
    'h8aa : romdata_int = 'h131d;
    'h8ab : romdata_int = 'h2721;
    'h8ac : romdata_int = 'h364d;
    'h8ad : romdata_int = 'h3639;
    'h8ae : romdata_int = 'h366e;
    'h8af : romdata_int = 'h550a;
    'h8b0 : romdata_int = 'h7600;
    'h8b1 : romdata_int = 'h9f30;
    'h8b2 : romdata_int = 'h848; // Line descriptor for 3_5
    'h8b3 : romdata_int = 'h364;
    'h8b4 : romdata_int = 'hc7c;
    'h8b5 : romdata_int = 'h283e;
    'h8b6 : romdata_int = 'h2b52;
    'h8b7 : romdata_int = 'h3d32;
    'h8b8 : romdata_int = 'h4622;
    'h8b9 : romdata_int = 'h7800;
    'h8ba : romdata_int = 'h7d15;
    'h8bb : romdata_int = 'hac5a;
    'h8bc : romdata_int = 'h4848; // Line descriptor for 3_5
    'h8bd : romdata_int = 'h2f0;
    'h8be : romdata_int = 'h316;
    'h8bf : romdata_int = 'h16b0;
    'h8c0 : romdata_int = 'h22cf;
    'h8c1 : romdata_int = 'h3231;
    'h8c2 : romdata_int = 'h411c;
    'h8c3 : romdata_int = 'h66b8;
    'h8c4 : romdata_int = 'h7a00;
    'h8c5 : romdata_int = 'h993b;
    'h8c6 : romdata_int = 'h848; // Line descriptor for 3_5
    'h8c7 : romdata_int = 'h2b;
    'h8c8 : romdata_int = 'h1d13;
    'h8c9 : romdata_int = 'h2030;
    'h8ca : romdata_int = 'h22d4;
    'h8cb : romdata_int = 'h391c;
    'h8cc : romdata_int = 'h4615;
    'h8cd : romdata_int = 'h6925;
    'h8ce : romdata_int = 'h7c00;
    'h8cf : romdata_int = 'h9860;
    'h8d0 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h8d1 : romdata_int = 'h1;
    'h8d2 : romdata_int = 'hcb5;
    'h8d3 : romdata_int = 'h14cf;
    'h8d4 : romdata_int = 'h20b5;
    'h8d5 : romdata_int = 'h4033;
    'h8d6 : romdata_int = 'h4632;
    'h8d7 : romdata_int = 'h5698;
    'h8d8 : romdata_int = 'h7e00;
    'h8d9 : romdata_int = 'ha6d3;
    'h8da : romdata_int = 'h848; // Line descriptor for 3_5
    'h8db : romdata_int = 'h44c;
    'h8dc : romdata_int = 'h1440;
    'h8dd : romdata_int = 'h14ab;
    'h8de : romdata_int = 'h2485;
    'h8df : romdata_int = 'h3d3a;
    'h8e0 : romdata_int = 'h40fd;
    'h8e1 : romdata_int = 'h5e65;
    'h8e2 : romdata_int = 'h8000;
    'h8e3 : romdata_int = 'h915b;
    'h8e4 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h8e5 : romdata_int = 'h53d;
    'h8e6 : romdata_int = 'hb18;
    'h8e7 : romdata_int = 'h14e4;
    'h8e8 : romdata_int = 'h1737;
    'h8e9 : romdata_int = 'h365e;
    'h8ea : romdata_int = 'h3ce4;
    'h8eb : romdata_int = 'h7695;
    'h8ec : romdata_int = 'h8200;
    'h8ed : romdata_int = 'h9726;
    'h8ee : romdata_int = 'h848; // Line descriptor for 3_5
    'h8ef : romdata_int = 'h137;
    'h8f0 : romdata_int = 'h1049;
    'h8f1 : romdata_int = 'h10f1;
    'h8f2 : romdata_int = 'h1acb;
    'h8f3 : romdata_int = 'h2d61;
    'h8f4 : romdata_int = 'h3b49;
    'h8f5 : romdata_int = 'h6b3c;
    'h8f6 : romdata_int = 'h8400;
    'h8f7 : romdata_int = 'hc633;
    'h8f8 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h8f9 : romdata_int = 'h35c;
    'h8fa : romdata_int = 'h89a;
    'h8fb : romdata_int = 'h1480;
    'h8fc : romdata_int = 'h3517;
    'h8fd : romdata_int = 'h404b;
    'h8fe : romdata_int = 'h4296;
    'h8ff : romdata_int = 'h6854;
    'h900 : romdata_int = 'h8600;
    'h901 : romdata_int = 'haac7;
    'h902 : romdata_int = 'h848; // Line descriptor for 3_5
    'h903 : romdata_int = 'hd22;
    'h904 : romdata_int = 'hec5;
    'h905 : romdata_int = 'h2a13;
    'h906 : romdata_int = 'h2c87;
    'h907 : romdata_int = 'h2e8e;
    'h908 : romdata_int = 'h40df;
    'h909 : romdata_int = 'h84bc;
    'h90a : romdata_int = 'h8800;
    'h90b : romdata_int = 'hb07a;
    'h90c : romdata_int = 'h4848; // Line descriptor for 3_5
    'h90d : romdata_int = 'h499;
    'h90e : romdata_int = 'h747;
    'h90f : romdata_int = 'h10c1;
    'h910 : romdata_int = 'h1d4d;
    'h911 : romdata_int = 'h2155;
    'h912 : romdata_int = 'h3d4f;
    'h913 : romdata_int = 'h4c95;
    'h914 : romdata_int = 'h8a00;
    'h915 : romdata_int = 'ha69c;
    'h916 : romdata_int = 'h848; // Line descriptor for 3_5
    'h917 : romdata_int = 'ha1;
    'h918 : romdata_int = 'h648;
    'h919 : romdata_int = 'hc5e;
    'h91a : romdata_int = 'h26b8;
    'h91b : romdata_int = 'h2e52;
    'h91c : romdata_int = 'h2eee;
    'h91d : romdata_int = 'h5707;
    'h91e : romdata_int = 'h8c00;
    'h91f : romdata_int = 'hc873;
    'h920 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h921 : romdata_int = 'h2;
    'h922 : romdata_int = 'h6a0;
    'h923 : romdata_int = 'h6ae;
    'h924 : romdata_int = 'h1aa4;
    'h925 : romdata_int = 'h314b;
    'h926 : romdata_int = 'h3744;
    'h927 : romdata_int = 'h4901;
    'h928 : romdata_int = 'h8e00;
    'h929 : romdata_int = 'hc0f1;
    'h92a : romdata_int = 'h848; // Line descriptor for 3_5
    'h92b : romdata_int = 'h20b;
    'h92c : romdata_int = 'h80f;
    'h92d : romdata_int = 'ha5a;
    'h92e : romdata_int = 'h1a0a;
    'h92f : romdata_int = 'h3029;
    'h930 : romdata_int = 'h3525;
    'h931 : romdata_int = 'h5f33;
    'h932 : romdata_int = 'h9000;
    'h933 : romdata_int = 'hd431;
    'h934 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h935 : romdata_int = 'h2a1;
    'h936 : romdata_int = 'had0;
    'h937 : romdata_int = 'h2067;
    'h938 : romdata_int = 'h234f;
    'h939 : romdata_int = 'h26ef;
    'h93a : romdata_int = 'h3065;
    'h93b : romdata_int = 'h823b;
    'h93c : romdata_int = 'h9200;
    'h93d : romdata_int = 'hcf13;
    'h93e : romdata_int = 'h848; // Line descriptor for 3_5
    'h93f : romdata_int = 'h133f;
    'h940 : romdata_int = 'h16fd;
    'h941 : romdata_int = 'h1915;
    'h942 : romdata_int = 'h3344;
    'h943 : romdata_int = 'h450a;
    'h944 : romdata_int = 'h46c0;
    'h945 : romdata_int = 'h5915;
    'h946 : romdata_int = 'h9400;
    'h947 : romdata_int = 'h9444;
    'h948 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h949 : romdata_int = 'h1e67;
    'h94a : romdata_int = 'h28e4;
    'h94b : romdata_int = 'h292f;
    'h94c : romdata_int = 'h2c77;
    'h94d : romdata_int = 'h3a7b;
    'h94e : romdata_int = 'h3c37;
    'h94f : romdata_int = 'h5520;
    'h950 : romdata_int = 'h9600;
    'h951 : romdata_int = 'hac21;
    'h952 : romdata_int = 'h848; // Line descriptor for 3_5
    'h953 : romdata_int = 'h166b;
    'h954 : romdata_int = 'h1e0f;
    'h955 : romdata_int = 'h28d5;
    'h956 : romdata_int = 'h2962;
    'h957 : romdata_int = 'h3215;
    'h958 : romdata_int = 'h3462;
    'h959 : romdata_int = 'h752e;
    'h95a : romdata_int = 'h9800;
    'h95b : romdata_int = 'hd0a8;
    'h95c : romdata_int = 'h4848; // Line descriptor for 3_5
    'h95d : romdata_int = 'h8e5;
    'h95e : romdata_int = 'h1228;
    'h95f : romdata_int = 'h330b;
    'h960 : romdata_int = 'h3355;
    'h961 : romdata_int = 'h3c48;
    'h962 : romdata_int = 'h455a;
    'h963 : romdata_int = 'h629a;
    'h964 : romdata_int = 'h9a00;
    'h965 : romdata_int = 'hbabb;
    'h966 : romdata_int = 'h848; // Line descriptor for 3_5
    'h967 : romdata_int = 'h28;
    'h968 : romdata_int = 'h49d;
    'h969 : romdata_int = 'h1418;
    'h96a : romdata_int = 'h2d47;
    'h96b : romdata_int = 'h3a8a;
    'h96c : romdata_int = 'h3f20;
    'h96d : romdata_int = 'h50b9;
    'h96e : romdata_int = 'h9c00;
    'h96f : romdata_int = 'ha351;
    'h970 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h971 : romdata_int = 'h8c4;
    'h972 : romdata_int = 'h1810;
    'h973 : romdata_int = 'h2470;
    'h974 : romdata_int = 'h30b5;
    'h975 : romdata_int = 'h4420;
    'h976 : romdata_int = 'h449c;
    'h977 : romdata_int = 'h8b10;
    'h978 : romdata_int = 'h9e00;
    'h979 : romdata_int = 'hb0c8;
    'h97a : romdata_int = 'h848; // Line descriptor for 3_5
    'h97b : romdata_int = 'h1037;
    'h97c : romdata_int = 'h112a;
    'h97d : romdata_int = 'h18ad;
    'h97e : romdata_int = 'h1f5e;
    'h97f : romdata_int = 'h28c7;
    'h980 : romdata_int = 'h3511;
    'h981 : romdata_int = 'h8084;
    'h982 : romdata_int = 'ha000;
    'h983 : romdata_int = 'ha4c2;
    'h984 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h985 : romdata_int = 'h42a;
    'h986 : romdata_int = 'h124e;
    'h987 : romdata_int = 'h2557;
    'h988 : romdata_int = 'h3c6b;
    'h989 : romdata_int = 'h3d37;
    'h98a : romdata_int = 'h4276;
    'h98b : romdata_int = 'h6f0d;
    'h98c : romdata_int = 'ha200;
    'h98d : romdata_int = 'hd428;
    'h98e : romdata_int = 'h848; // Line descriptor for 3_5
    'h98f : romdata_int = 'h101e;
    'h990 : romdata_int = 'h1158;
    'h991 : romdata_int = 'h30b6;
    'h992 : romdata_int = 'h314c;
    'h993 : romdata_int = 'h4259;
    'h994 : romdata_int = 'h4463;
    'h995 : romdata_int = 'h82f3;
    'h996 : romdata_int = 'h9a68;
    'h997 : romdata_int = 'ha400;
    'h998 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h999 : romdata_int = 'he7d;
    'h99a : romdata_int = 'h1a32;
    'h99b : romdata_int = 'h2b44;
    'h99c : romdata_int = 'h344e;
    'h99d : romdata_int = 'h3505;
    'h99e : romdata_int = 'h4627;
    'h99f : romdata_int = 'h6d12;
    'h9a0 : romdata_int = 'ha600;
    'h9a1 : romdata_int = 'hb638;
    'h9a2 : romdata_int = 'h848; // Line descriptor for 3_5
    'h9a3 : romdata_int = 'h923;
    'h9a4 : romdata_int = 'h1906;
    'h9a5 : romdata_int = 'h1b3e;
    'h9a6 : romdata_int = 'h2ab3;
    'h9a7 : romdata_int = 'h2b62;
    'h9a8 : romdata_int = 'h3736;
    'h9a9 : romdata_int = 'h8ef0;
    'h9aa : romdata_int = 'h90c1;
    'h9ab : romdata_int = 'ha800;
    'h9ac : romdata_int = 'h4848; // Line descriptor for 3_5
    'h9ad : romdata_int = 'h734;
    'h9ae : romdata_int = 'h1312;
    'h9af : romdata_int = 'h1ab3;
    'h9b0 : romdata_int = 'h2818;
    'h9b1 : romdata_int = 'h2ef7;
    'h9b2 : romdata_int = 'h3838;
    'h9b3 : romdata_int = 'h7032;
    'h9b4 : romdata_int = 'h9338;
    'h9b5 : romdata_int = 'haa00;
    'h9b6 : romdata_int = 'h848; // Line descriptor for 3_5
    'h9b7 : romdata_int = 'ha83;
    'h9b8 : romdata_int = 'hee9;
    'h9b9 : romdata_int = 'h1c0b;
    'h9ba : romdata_int = 'h28fc;
    'h9bb : romdata_int = 'h3b47;
    'h9bc : romdata_int = 'h4089;
    'h9bd : romdata_int = 'h4a29;
    'h9be : romdata_int = 'hac00;
    'h9bf : romdata_int = 'hd62f;
    'h9c0 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h9c1 : romdata_int = 'h338;
    'h9c2 : romdata_int = 'h1916;
    'h9c3 : romdata_int = 'h1c45;
    'h9c4 : romdata_int = 'h2e4b;
    'h9c5 : romdata_int = 'h4308;
    'h9c6 : romdata_int = 'h4558;
    'h9c7 : romdata_int = 'h72b9;
    'h9c8 : romdata_int = 'ha8d7;
    'h9c9 : romdata_int = 'hae00;
    'h9ca : romdata_int = 'h848; // Line descriptor for 3_5
    'h9cb : romdata_int = 'he4c;
    'h9cc : romdata_int = 'h1c7a;
    'h9cd : romdata_int = 'h2a38;
    'h9ce : romdata_int = 'h2a75;
    'h9cf : romdata_int = 'h2edf;
    'h9d0 : romdata_int = 'h4291;
    'h9d1 : romdata_int = 'h4e6c;
    'h9d2 : romdata_int = 'haf5a;
    'h9d3 : romdata_int = 'hb000;
    'h9d4 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h9d5 : romdata_int = 'h115;
    'h9d6 : romdata_int = 'hf4a;
    'h9d7 : romdata_int = 'h1221;
    'h9d8 : romdata_int = 'h1338;
    'h9d9 : romdata_int = 'h1a72;
    'h9da : romdata_int = 'h3844;
    'h9db : romdata_int = 'h7a33;
    'h9dc : romdata_int = 'h9cb1;
    'h9dd : romdata_int = 'hb200;
    'h9de : romdata_int = 'h848; // Line descriptor for 3_5
    'h9df : romdata_int = 'h20cb;
    'h9e0 : romdata_int = 'h2080;
    'h9e1 : romdata_int = 'h20e5;
    'h9e2 : romdata_int = 'h2233;
    'h9e3 : romdata_int = 'h275f;
    'h9e4 : romdata_int = 'h4023;
    'h9e5 : romdata_int = 'h8942;
    'h9e6 : romdata_int = 'hb400;
    'h9e7 : romdata_int = 'hd26b;
    'h9e8 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h9e9 : romdata_int = 'h259;
    'h9ea : romdata_int = 'h1923;
    'h9eb : romdata_int = 'h24e6;
    'h9ec : romdata_int = 'h366f;
    'h9ed : romdata_int = 'h3ab7;
    'h9ee : romdata_int = 'h3ea4;
    'h9ef : romdata_int = 'h7e4f;
    'h9f0 : romdata_int = 'hb600;
    'h9f1 : romdata_int = 'hcb16;
    'h9f2 : romdata_int = 'h848; // Line descriptor for 3_5
    'h9f3 : romdata_int = 'h1e41;
    'h9f4 : romdata_int = 'h2032;
    'h9f5 : romdata_int = 'h2559;
    'h9f6 : romdata_int = 'h2567;
    'h9f7 : romdata_int = 'h2c01;
    'h9f8 : romdata_int = 'h2c19;
    'h9f9 : romdata_int = 'h88a1;
    'h9fa : romdata_int = 'hb800;
    'h9fb : romdata_int = 'hd33c;
    'h9fc : romdata_int = 'h4848; // Line descriptor for 3_5
    'h9fd : romdata_int = 'h4ef;
    'h9fe : romdata_int = 'h1308;
    'h9ff : romdata_int = 'h1855;
    'ha00 : romdata_int = 'h20db;
    'ha01 : romdata_int = 'h2633;
    'ha02 : romdata_int = 'h4464;
    'ha03 : romdata_int = 'h7a58;
    'ha04 : romdata_int = 'haa82;
    'ha05 : romdata_int = 'hba00;
    'ha06 : romdata_int = 'h848; // Line descriptor for 3_5
    'ha07 : romdata_int = 'h8e;
    'ha08 : romdata_int = 'ha0e;
    'ha09 : romdata_int = 'h32f4;
    'ha0a : romdata_int = 'h3864;
    'ha0b : romdata_int = 'h3e6e;
    'ha0c : romdata_int = 'h4428;
    'ha0d : romdata_int = 'h8618;
    'ha0e : romdata_int = 'hbc00;
    'ha0f : romdata_int = 'hbe15;
    'ha10 : romdata_int = 'h4848; // Line descriptor for 3_5
    'ha11 : romdata_int = 'h760;
    'ha12 : romdata_int = 'h894;
    'ha13 : romdata_int = 'hac5;
    'ha14 : romdata_int = 'h194c;
    'ha15 : romdata_int = 'h2149;
    'ha16 : romdata_int = 'h2646;
    'ha17 : romdata_int = 'h4eaa;
    'ha18 : romdata_int = 'h94ae;
    'ha19 : romdata_int = 'hbe00;
    'ha1a : romdata_int = 'h848; // Line descriptor for 3_5
    'ha1b : romdata_int = 'h4c7;
    'ha1c : romdata_int = 'hd34;
    'ha1d : romdata_int = 'h32fa;
    'ha1e : romdata_int = 'h3861;
    'ha1f : romdata_int = 'h429e;
    'ha20 : romdata_int = 'h46d0;
    'ha21 : romdata_int = 'h8ebe;
    'ha22 : romdata_int = 'ha00f;
    'ha23 : romdata_int = 'hc000;
    'ha24 : romdata_int = 'h4848; // Line descriptor for 3_5
    'ha25 : romdata_int = 'h711;
    'ha26 : romdata_int = 'hae7;
    'ha27 : romdata_int = 'h1d51;
    'ha28 : romdata_int = 'h251a;
    'ha29 : romdata_int = 'h28ad;
    'ha2a : romdata_int = 'h2b35;
    'ha2b : romdata_int = 'h64bf;
    'ha2c : romdata_int = 'hc200;
    'ha2d : romdata_int = 'hc812;
    'ha2e : romdata_int = 'h848; // Line descriptor for 3_5
    'ha2f : romdata_int = 'h72;
    'ha30 : romdata_int = 'h183c;
    'ha31 : romdata_int = 'h3b28;
    'ha32 : romdata_int = 'h3cb8;
    'ha33 : romdata_int = 'h409c;
    'ha34 : romdata_int = 'h42e3;
    'ha35 : romdata_int = 'h4a91;
    'ha36 : romdata_int = 'ha840;
    'ha37 : romdata_int = 'hc400;
    'ha38 : romdata_int = 'h4848; // Line descriptor for 3_5
    'ha39 : romdata_int = 'h339;
    'ha3a : romdata_int = 'h84e;
    'ha3b : romdata_int = 'h2d5c;
    'ha3c : romdata_int = 'h3953;
    'ha3d : romdata_int = 'h3f65;
    'ha3e : romdata_int = 'h413c;
    'ha3f : romdata_int = 'h8539;
    'ha40 : romdata_int = 'h925c;
    'ha41 : romdata_int = 'hc600;
    'ha42 : romdata_int = 'h848; // Line descriptor for 3_5
    'ha43 : romdata_int = 'hc5f;
    'ha44 : romdata_int = 'h10e5;
    'ha45 : romdata_int = 'h1498;
    'ha46 : romdata_int = 'h2f25;
    'ha47 : romdata_int = 'h44e1;
    'ha48 : romdata_int = 'h4741;
    'ha49 : romdata_int = 'h5a9c;
    'ha4a : romdata_int = 'h9d52;
    'ha4b : romdata_int = 'hc800;
    'ha4c : romdata_int = 'h4848; // Line descriptor for 3_5
    'ha4d : romdata_int = 'hf11;
    'ha4e : romdata_int = 'h1c99;
    'ha4f : romdata_int = 'h22eb;
    'ha50 : romdata_int = 'h34c2;
    'ha51 : romdata_int = 'h3eec;
    'ha52 : romdata_int = 'h4652;
    'ha53 : romdata_int = 'h8cbc;
    'ha54 : romdata_int = 'hca00;
    'ha55 : romdata_int = 'hd66b;
    'ha56 : romdata_int = 'h848; // Line descriptor for 3_5
    'ha57 : romdata_int = 'ha13;
    'ha58 : romdata_int = 'h2755;
    'ha59 : romdata_int = 'h28f2;
    'ha5a : romdata_int = 'h2a58;
    'ha5b : romdata_int = 'h3154;
    'ha5c : romdata_int = 'h3ac4;
    'ha5d : romdata_int = 'h8cba;
    'ha5e : romdata_int = 'haf56;
    'ha5f : romdata_int = 'hcc00;
    'ha60 : romdata_int = 'h4848; // Line descriptor for 3_5
    'ha61 : romdata_int = 'hcd9;
    'ha62 : romdata_int = 'hd2b;
    'ha63 : romdata_int = 'h1425;
    'ha64 : romdata_int = 'h3893;
    'ha65 : romdata_int = 'h424f;
    'ha66 : romdata_int = 'h44af;
    'ha67 : romdata_int = 'h5d1e;
    'ha68 : romdata_int = 'hb211;
    'ha69 : romdata_int = 'hce00;
    'ha6a : romdata_int = 'h848; // Line descriptor for 3_5
    'ha6b : romdata_int = 'h8d8;
    'ha6c : romdata_int = 'ha77;
    'ha6d : romdata_int = 'hc06;
    'ha6e : romdata_int = 'h1c6f;
    'ha6f : romdata_int = 'h233b;
    'ha70 : romdata_int = 'h34ad;
    'ha71 : romdata_int = 'h6a50;
    'ha72 : romdata_int = 'hbe53;
    'ha73 : romdata_int = 'hd000;
    'ha74 : romdata_int = 'h4848; // Line descriptor for 3_5
    'ha75 : romdata_int = 'h1761;
    'ha76 : romdata_int = 'h1958;
    'ha77 : romdata_int = 'h24ba;
    'ha78 : romdata_int = 'h271c;
    'ha79 : romdata_int = 'h38c6;
    'ha7a : romdata_int = 'h4607;
    'ha7b : romdata_int = 'h6131;
    'ha7c : romdata_int = 'hba54;
    'ha7d : romdata_int = 'hd200;
    'ha7e : romdata_int = 'h848; // Line descriptor for 3_5
    'ha7f : romdata_int = 'h1a9a;
    'ha80 : romdata_int = 'h2137;
    'ha81 : romdata_int = 'h2688;
    'ha82 : romdata_int = 'h3112;
    'ha83 : romdata_int = 'h380e;
    'ha84 : romdata_int = 'h383b;
    'ha85 : romdata_int = 'h5cd0;
    'ha86 : romdata_int = 'hb520;
    'ha87 : romdata_int = 'hd400;
    'ha88 : romdata_int = 'h6848; // Line descriptor for 3_5
    'ha89 : romdata_int = 'h140a;
    'ha8a : romdata_int = 'h1e4c;
    'ha8b : romdata_int = 'h26c4;
    'ha8c : romdata_int = 'h2a70;
    'ha8d : romdata_int = 'h2b21;
    'ha8e : romdata_int = 'h3f55;
    'ha8f : romdata_int = 'h6c3a;
    'ha90 : romdata_int = 'hc51d;
    'ha91 : romdata_int = 'hd600;
    'ha92 : romdata_int = 'h73c; // Line descriptor for 2_3
    'ha93 : romdata_int = 'h0;
    'ha94 : romdata_int = 'h4;
    'ha95 : romdata_int = 'h16ec;
    'ha96 : romdata_int = 'h18e6;
    'ha97 : romdata_int = 'h4f1c;
    'ha98 : romdata_int = 'h7800;
    'ha99 : romdata_int = 'h9ea5;
    'ha9a : romdata_int = 'h9ee8;
    'ha9b : romdata_int = 'h473c; // Line descriptor for 2_3
    'ha9c : romdata_int = 'h200;
    'ha9d : romdata_int = 'h6bd;
    'ha9e : romdata_int = 'hf37;
    'ha9f : romdata_int = 'h18ec;
    'haa0 : romdata_int = 'h22e1;
    'haa1 : romdata_int = 'h7a00;
    'haa2 : romdata_int = 'hde3d;
    'haa3 : romdata_int = 'he12e;
    'haa4 : romdata_int = 'h73c; // Line descriptor for 2_3
    'haa5 : romdata_int = 'h400;
    'haa6 : romdata_int = 'h1097;
    'haa7 : romdata_int = 'h1648;
    'haa8 : romdata_int = 'h4f3e;
    'haa9 : romdata_int = 'h5f5f;
    'haaa : romdata_int = 'h7c00;
    'haab : romdata_int = 'haa48;
    'haac : romdata_int = 'hea70;
    'haad : romdata_int = 'h473c; // Line descriptor for 2_3
    'haae : romdata_int = 'h334;
    'haaf : romdata_int = 'h600;
    'hab0 : romdata_int = 'h667;
    'hab1 : romdata_int = 'hce5;
    'hab2 : romdata_int = 'h2013;
    'hab3 : romdata_int = 'h7e00;
    'hab4 : romdata_int = 'hd50b;
    'hab5 : romdata_int = 'he52c;
    'hab6 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hab7 : romdata_int = 'h261;
    'hab8 : romdata_int = 'h4c9;
    'hab9 : romdata_int = 'h800;
    'haba : romdata_int = 'h3d53;
    'habb : romdata_int = 'h741f;
    'habc : romdata_int = 'h8000;
    'habd : romdata_int = 'h910a;
    'habe : romdata_int = 'h9c22;
    'habf : romdata_int = 'h473c; // Line descriptor for 2_3
    'hac0 : romdata_int = 'ha00;
    'hac1 : romdata_int = 'hb38;
    'hac2 : romdata_int = 'he5c;
    'hac3 : romdata_int = 'h129e;
    'hac4 : romdata_int = 'h72a4;
    'hac5 : romdata_int = 'h7c33;
    'hac6 : romdata_int = 'h8200;
    'hac7 : romdata_int = 'h84c1;
    'hac8 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hac9 : romdata_int = 'h89;
    'haca : romdata_int = 'hc00;
    'hacb : romdata_int = 'hc08;
    'hacc : romdata_int = 'h10d5;
    'hacd : romdata_int = 'h4660;
    'hace : romdata_int = 'h8400;
    'hacf : romdata_int = 'h8a14;
    'had0 : romdata_int = 'ha6a2;
    'had1 : romdata_int = 'h473c; // Line descriptor for 2_3
    'had2 : romdata_int = 'h2e;
    'had3 : romdata_int = 'h2e0;
    'had4 : romdata_int = 'he00;
    'had5 : romdata_int = 'hf58;
    'had6 : romdata_int = 'h1d0b;
    'had7 : romdata_int = 'h8600;
    'had8 : romdata_int = 'hb07b;
    'had9 : romdata_int = 'hc71e;
    'hada : romdata_int = 'h73c; // Line descriptor for 2_3
    'hadb : romdata_int = 'h1000;
    'hadc : romdata_int = 'h1406;
    'hadd : romdata_int = 'h16d2;
    'hade : romdata_int = 'h1a31;
    'hadf : romdata_int = 'h3ef3;
    'hae0 : romdata_int = 'h8800;
    'hae1 : romdata_int = 'hd654;
    'hae2 : romdata_int = 'hdd0d;
    'hae3 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hae4 : romdata_int = 'h948;
    'hae5 : romdata_int = 'hace;
    'hae6 : romdata_int = 'heb0;
    'hae7 : romdata_int = 'h1200;
    'hae8 : romdata_int = 'h5468;
    'hae9 : romdata_int = 'h8a00;
    'haea : romdata_int = 'hbc1a;
    'haeb : romdata_int = 'hcf33;
    'haec : romdata_int = 'h73c; // Line descriptor for 2_3
    'haed : romdata_int = 'hccf;
    'haee : romdata_int = 'he87;
    'haef : romdata_int = 'h1400;
    'haf0 : romdata_int = 'h4c44;
    'haf1 : romdata_int = 'h553d;
    'haf2 : romdata_int = 'h8c00;
    'haf3 : romdata_int = 'haa85;
    'haf4 : romdata_int = 'hbc7d;
    'haf5 : romdata_int = 'h473c; // Line descriptor for 2_3
    'haf6 : romdata_int = 'h477;
    'haf7 : romdata_int = 'hc5d;
    'haf8 : romdata_int = 'h103f;
    'haf9 : romdata_int = 'h1600;
    'hafa : romdata_int = 'h4344;
    'hafb : romdata_int = 'h8e00;
    'hafc : romdata_int = 'ha466;
    'hafd : romdata_int = 'hc203;
    'hafe : romdata_int = 'h73c; // Line descriptor for 2_3
    'haff : romdata_int = 'h6a6;
    'hb00 : romdata_int = 'h1351;
    'hb01 : romdata_int = 'h1800;
    'hb02 : romdata_int = 'h58c4;
    'hb03 : romdata_int = 'h7028;
    'hb04 : romdata_int = 'h7f30;
    'hb05 : romdata_int = 'h9000;
    'hb06 : romdata_int = 'hce8d;
    'hb07 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb08 : romdata_int = 'h137;
    'hb09 : romdata_int = 'h26b;
    'hb0a : romdata_int = 'h1643;
    'hb0b : romdata_int = 'h1a00;
    'hb0c : romdata_int = 'h5151;
    'hb0d : romdata_int = 'h82a9;
    'hb0e : romdata_int = 'h9200;
    'hb0f : romdata_int = 'h9804;
    'hb10 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hb11 : romdata_int = 'h4d5;
    'hb12 : romdata_int = 'h92a;
    'hb13 : romdata_int = 'h1c00;
    'hb14 : romdata_int = 'h2ed2;
    'hb15 : romdata_int = 'h3711;
    'hb16 : romdata_int = 'h9400;
    'hb17 : romdata_int = 'h9a15;
    'hb18 : romdata_int = 'ha45a;
    'hb19 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb1a : romdata_int = 'h44a;
    'hb1b : romdata_int = 'h140f;
    'hb1c : romdata_int = 'h1e00;
    'hb1d : romdata_int = 'h3325;
    'hb1e : romdata_int = 'h7120;
    'hb1f : romdata_int = 'h8e9c;
    'hb20 : romdata_int = 'h9600;
    'hb21 : romdata_int = 'hd725;
    'hb22 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hb23 : romdata_int = 'h6f2;
    'hb24 : romdata_int = 'h14e2;
    'hb25 : romdata_int = 'h2000;
    'hb26 : romdata_int = 'h2767;
    'hb27 : romdata_int = 'h4408;
    'hb28 : romdata_int = 'h9800;
    'hb29 : romdata_int = 'had04;
    'hb2a : romdata_int = 'hcc54;
    'hb2b : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb2c : romdata_int = 'h52b;
    'hb2d : romdata_int = 'ha21;
    'hb2e : romdata_int = 'hcc0;
    'hb2f : romdata_int = 'h2200;
    'hb30 : romdata_int = 'h4446;
    'hb31 : romdata_int = 'h9a00;
    'hb32 : romdata_int = 'h9cf6;
    'hb33 : romdata_int = 'hd850;
    'hb34 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hb35 : romdata_int = 'hafd;
    'hb36 : romdata_int = 'h1313;
    'hb37 : romdata_int = 'h2400;
    'hb38 : romdata_int = 'h3a6f;
    'hb39 : romdata_int = 'h4c61;
    'hb3a : romdata_int = 'h8497;
    'hb3b : romdata_int = 'h9c00;
    'hb3c : romdata_int = 'hb159;
    'hb3d : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb3e : romdata_int = 'hb0;
    'hb3f : romdata_int = 'h134d;
    'hb40 : romdata_int = 'h2600;
    'hb41 : romdata_int = 'h5ec4;
    'hb42 : romdata_int = 'h6437;
    'hb43 : romdata_int = 'h8659;
    'hb44 : romdata_int = 'h9e00;
    'hb45 : romdata_int = 'ha85b;
    'hb46 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hb47 : romdata_int = 'h255;
    'hb48 : romdata_int = 'ha1c;
    'hb49 : romdata_int = 'h2096;
    'hb4a : romdata_int = 'h2800;
    'hb4b : romdata_int = 'h5949;
    'hb4c : romdata_int = 'h7a9c;
    'hb4d : romdata_int = 'ha000;
    'hb4e : romdata_int = 'hb42b;
    'hb4f : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb50 : romdata_int = 'heca;
    'hb51 : romdata_int = 'hf33;
    'hb52 : romdata_int = 'h2a00;
    'hb53 : romdata_int = 'h3874;
    'hb54 : romdata_int = 'h48af;
    'hb55 : romdata_int = 'ha200;
    'hb56 : romdata_int = 'ha2a5;
    'hb57 : romdata_int = 'haf03;
    'hb58 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hb59 : romdata_int = 'h688;
    'hb5a : romdata_int = 'h10a1;
    'hb5b : romdata_int = 'h2c00;
    'hb5c : romdata_int = 'h60a1;
    'hb5d : romdata_int = 'h6e56;
    'hb5e : romdata_int = 'h8c12;
    'hb5f : romdata_int = 'h9485;
    'hb60 : romdata_int = 'ha400;
    'hb61 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb62 : romdata_int = 'h10b;
    'hb63 : romdata_int = 'h866;
    'hb64 : romdata_int = 'h16aa;
    'hb65 : romdata_int = 'h2e00;
    'hb66 : romdata_int = 'h6a63;
    'hb67 : romdata_int = 'ha600;
    'hb68 : romdata_int = 'he633;
    'hb69 : romdata_int = 'he658;
    'hb6a : romdata_int = 'h73c; // Line descriptor for 2_3
    'hb6b : romdata_int = 'h464;
    'hb6c : romdata_int = 'h10fe;
    'hb6d : romdata_int = 'h1766;
    'hb6e : romdata_int = 'h3000;
    'hb6f : romdata_int = 'h5b47;
    'hb70 : romdata_int = 'h8896;
    'hb71 : romdata_int = 'ha800;
    'hb72 : romdata_int = 'hb339;
    'hb73 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb74 : romdata_int = 'h86;
    'hb75 : romdata_int = 'h2e6;
    'hb76 : romdata_int = 'h1345;
    'hb77 : romdata_int = 'h3200;
    'hb78 : romdata_int = 'h4ac6;
    'hb79 : romdata_int = 'haa00;
    'hb7a : romdata_int = 'hc537;
    'hb7b : romdata_int = 'hd310;
    'hb7c : romdata_int = 'h73c; // Line descriptor for 2_3
    'hb7d : romdata_int = 'h8;
    'hb7e : romdata_int = 'h858;
    'hb7f : romdata_int = 'h3400;
    'hb80 : romdata_int = 'h6c7a;
    'hb81 : romdata_int = 'h6cc3;
    'hb82 : romdata_int = 'h9b41;
    'hb83 : romdata_int = 'ha32f;
    'hb84 : romdata_int = 'hac00;
    'hb85 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb86 : romdata_int = 'h31e;
    'hb87 : romdata_int = 'h916;
    'hb88 : romdata_int = 'h3600;
    'hb89 : romdata_int = 'h3cd8;
    'hb8a : romdata_int = 'h746f;
    'hb8b : romdata_int = 'h9064;
    'hb8c : romdata_int = 'hae00;
    'hb8d : romdata_int = 'hc098;
    'hb8e : romdata_int = 'h73c; // Line descriptor for 2_3
    'hb8f : romdata_int = 'h536;
    'hb90 : romdata_int = 'h143a;
    'hb91 : romdata_int = 'h144c;
    'hb92 : romdata_int = 'h2ca7;
    'hb93 : romdata_int = 'h3800;
    'hb94 : romdata_int = 'hb000;
    'hb95 : romdata_int = 'hd2d4;
    'hb96 : romdata_int = 'he295;
    'hb97 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb98 : romdata_int = 'h1299;
    'hb99 : romdata_int = 'h1689;
    'hb9a : romdata_int = 'h387b;
    'hb9b : romdata_int = 'h3a00;
    'hb9c : romdata_int = 'h6e5d;
    'hb9d : romdata_int = 'h92f6;
    'hb9e : romdata_int = 'hb200;
    'hb9f : romdata_int = 'hb72a;
    'hba0 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hba1 : romdata_int = 'hb19;
    'hba2 : romdata_int = 'h126f;
    'hba3 : romdata_int = 'h2424;
    'hba4 : romdata_int = 'h3c00;
    'hba5 : romdata_int = 'h4679;
    'hba6 : romdata_int = 'hac5c;
    'hba7 : romdata_int = 'hb400;
    'hba8 : romdata_int = 'hc315;
    'hba9 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hbaa : romdata_int = 'h84d;
    'hbab : romdata_int = 'hd22;
    'hbac : romdata_int = 'heee;
    'hbad : romdata_int = 'h160a;
    'hbae : romdata_int = 'h3e00;
    'hbaf : romdata_int = 'hb600;
    'hbb0 : romdata_int = 'hc838;
    'hbb1 : romdata_int = 'hea4f;
    'hbb2 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hbb3 : romdata_int = 'h2d5;
    'hbb4 : romdata_int = 'ha2a;
    'hbb5 : romdata_int = 'he88;
    'hbb6 : romdata_int = 'h16ea;
    'hbb7 : romdata_int = 'h4000;
    'hbb8 : romdata_int = 'h926b;
    'hbb9 : romdata_int = 'ha007;
    'hbba : romdata_int = 'hb800;
    'hbbb : romdata_int = 'h473c; // Line descriptor for 2_3
    'hbbc : romdata_int = 'h28a;
    'hbbd : romdata_int = 'h127a;
    'hbbe : romdata_int = 'h14b8;
    'hbbf : romdata_int = 'h3462;
    'hbc0 : romdata_int = 'h4200;
    'hbc1 : romdata_int = 'hba00;
    'hbc2 : romdata_int = 'hd0c9;
    'hbc3 : romdata_int = 'he2c4;
    'hbc4 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hbc5 : romdata_int = 'h722;
    'hbc6 : romdata_int = 'hec3;
    'hbc7 : romdata_int = 'h4400;
    'hbc8 : romdata_int = 'h6883;
    'hbc9 : romdata_int = 'h7355;
    'hbca : romdata_int = 'h82b2;
    'hbcb : romdata_int = 'h8b10;
    'hbcc : romdata_int = 'hbc00;
    'hbcd : romdata_int = 'h473c; // Line descriptor for 2_3
    'hbce : romdata_int = 'h462;
    'hbcf : romdata_int = 'h16ce;
    'hbd0 : romdata_int = 'h2e08;
    'hbd1 : romdata_int = 'h348d;
    'hbd2 : romdata_int = 'h4600;
    'hbd3 : romdata_int = 'h889e;
    'hbd4 : romdata_int = 'hbe00;
    'hbd5 : romdata_int = 'hd93c;
    'hbd6 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hbd7 : romdata_int = 'h65c;
    'hbd8 : romdata_int = 'hac9;
    'hbd9 : romdata_int = 'h26cb;
    'hbda : romdata_int = 'h4800;
    'hbdb : romdata_int = 'h6648;
    'hbdc : romdata_int = 'h8f5a;
    'hbdd : romdata_int = 'hb66c;
    'hbde : romdata_int = 'hc000;
    'hbdf : romdata_int = 'h473c; // Line descriptor for 2_3
    'hbe0 : romdata_int = 'h554;
    'hbe1 : romdata_int = 'h749;
    'hbe2 : romdata_int = 'h1281;
    'hbe3 : romdata_int = 'h294b;
    'hbe4 : romdata_int = 'h4a00;
    'hbe5 : romdata_int = 'hc200;
    'hbe6 : romdata_int = 'hc503;
    'hbe7 : romdata_int = 'hc75c;
    'hbe8 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hbe9 : romdata_int = 'h8f3;
    'hbea : romdata_int = 'h128b;
    'hbeb : romdata_int = 'h2a84;
    'hbec : romdata_int = 'h412a;
    'hbed : romdata_int = 'h4c00;
    'hbee : romdata_int = 'hb801;
    'hbef : romdata_int = 'hc400;
    'hbf0 : romdata_int = 'hcc99;
    'hbf1 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hbf2 : romdata_int = 'h9a;
    'hbf3 : romdata_int = 'h174c;
    'hbf4 : romdata_int = 'h3b09;
    'hbf5 : romdata_int = 'h4b53;
    'hbf6 : romdata_int = 'h4e00;
    'hbf7 : romdata_int = 'hbb56;
    'hbf8 : romdata_int = 'hc600;
    'hbf9 : romdata_int = 'hde32;
    'hbfa : romdata_int = 'h73c; // Line descriptor for 2_3
    'hbfb : romdata_int = 'h2a5;
    'hbfc : romdata_int = 'he45;
    'hbfd : romdata_int = 'h2d09;
    'hbfe : romdata_int = 'h5000;
    'hbff : romdata_int = 'h6a48;
    'hc00 : romdata_int = 'hbf0a;
    'hc01 : romdata_int = 'hc800;
    'hc02 : romdata_int = 'hec84;
    'hc03 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc04 : romdata_int = 'h490;
    'hc05 : romdata_int = 'hf06;
    'hc06 : romdata_int = 'h308d;
    'hc07 : romdata_int = 'h5200;
    'hc08 : romdata_int = 'h5c3a;
    'hc09 : romdata_int = 'h8098;
    'hc0a : romdata_int = 'haeb1;
    'hc0b : romdata_int = 'hca00;
    'hc0c : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc0d : romdata_int = 'hb08;
    'hc0e : romdata_int = 'h1550;
    'hc0f : romdata_int = 'h1eb8;
    'hc10 : romdata_int = 'h5400;
    'hc11 : romdata_int = 'h60d9;
    'hc12 : romdata_int = 'h8104;
    'hc13 : romdata_int = 'h96f5;
    'hc14 : romdata_int = 'hcc00;
    'hc15 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc16 : romdata_int = 'hc18;
    'hc17 : romdata_int = 'h1234;
    'hc18 : romdata_int = 'h36ad;
    'hc19 : romdata_int = 'h426f;
    'hc1a : romdata_int = 'h5600;
    'hc1b : romdata_int = 'hc0ab;
    'hc1c : romdata_int = 'hce00;
    'hc1d : romdata_int = 'hdb12;
    'hc1e : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc1f : romdata_int = 'h267;
    'hc20 : romdata_int = 'h958;
    'hc21 : romdata_int = 'h3317;
    'hc22 : romdata_int = 'h5800;
    'hc23 : romdata_int = 'h7756;
    'hc24 : romdata_int = 'hb495;
    'hc25 : romdata_int = 'hba3d;
    'hc26 : romdata_int = 'hd000;
    'hc27 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc28 : romdata_int = 'hceb;
    'hc29 : romdata_int = 'h14b5;
    'hc2a : romdata_int = 'h4894;
    'hc2b : romdata_int = 'h5342;
    'hc2c : romdata_int = 'h5a00;
    'hc2d : romdata_int = 'h9832;
    'hc2e : romdata_int = 'ha8c8;
    'hc2f : romdata_int = 'hd200;
    'hc30 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc31 : romdata_int = 'hd5;
    'hc32 : romdata_int = 'h1140;
    'hc33 : romdata_int = 'h1f55;
    'hc34 : romdata_int = 'h5345;
    'hc35 : romdata_int = 'h5c00;
    'hc36 : romdata_int = 'h792f;
    'hc37 : romdata_int = 'h7a89;
    'hc38 : romdata_int = 'hd400;
    'hc39 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc3a : romdata_int = 'hc40;
    'hc3b : romdata_int = 'hcfd;
    'hc3c : romdata_int = 'h1aa0;
    'hc3d : romdata_int = 'h5e00;
    'hc3e : romdata_int = 'h64b8;
    'hc3f : romdata_int = 'h791e;
    'hc40 : romdata_int = 'hd600;
    'hc41 : romdata_int = 'he4df;
    'hc42 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc43 : romdata_int = 'h15c;
    'hc44 : romdata_int = 'h81a;
    'hc45 : romdata_int = 'h2419;
    'hc46 : romdata_int = 'h5a7b;
    'hc47 : romdata_int = 'h6000;
    'hc48 : romdata_int = 'hb8b9;
    'hc49 : romdata_int = 'hd800;
    'hc4a : romdata_int = 'he915;
    'hc4b : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc4c : romdata_int = 'h727;
    'hc4d : romdata_int = 'ha33;
    'hc4e : romdata_int = 'h146f;
    'hc4f : romdata_int = 'h2a45;
    'hc50 : romdata_int = 'h6200;
    'hc51 : romdata_int = 'h96ea;
    'hc52 : romdata_int = 'hda00;
    'hc53 : romdata_int = 'hee3b;
    'hc54 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc55 : romdata_int = 'h4b6;
    'hc56 : romdata_int = 'h10a6;
    'hc57 : romdata_int = 'h308c;
    'hc58 : romdata_int = 'h3e29;
    'hc59 : romdata_int = 'h6400;
    'hc5a : romdata_int = 'hdc00;
    'hc5b : romdata_int = 'he13c;
    'hc5c : romdata_int = 'heef3;
    'hc5d : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc5e : romdata_int = 'hae;
    'hc5f : romdata_int = 'ha50;
    'hc60 : romdata_int = 'hc65;
    'hc61 : romdata_int = 'h1560;
    'hc62 : romdata_int = 'h6600;
    'hc63 : romdata_int = 'h9535;
    'hc64 : romdata_int = 'hde00;
    'hc65 : romdata_int = 'he808;
    'hc66 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc67 : romdata_int = 'h734;
    'hc68 : romdata_int = 'h10a8;
    'hc69 : romdata_int = 'h50cd;
    'hc6a : romdata_int = 'h673a;
    'hc6b : romdata_int = 'h6800;
    'hc6c : romdata_int = 'hbec2;
    'hc6d : romdata_int = 'hcb4e;
    'hc6e : romdata_int = 'he000;
    'hc6f : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc70 : romdata_int = 'hc7b;
    'hc71 : romdata_int = 'h1511;
    'hc72 : romdata_int = 'h1cf4;
    'hc73 : romdata_int = 'h573f;
    'hc74 : romdata_int = 'h6a00;
    'hc75 : romdata_int = 'h7c75;
    'hc76 : romdata_int = 'hd159;
    'hc77 : romdata_int = 'he200;
    'hc78 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc79 : romdata_int = 'h105a;
    'hc7a : romdata_int = 'h1744;
    'hc7b : romdata_int = 'h2242;
    'hc7c : romdata_int = 'h6294;
    'hc7d : romdata_int = 'h6c00;
    'hc7e : romdata_int = 'h8cf9;
    'hc7f : romdata_int = 'ha07a;
    'hc80 : romdata_int = 'he400;
    'hc81 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc82 : romdata_int = 'h8ee;
    'hc83 : romdata_int = 'h10b1;
    'hc84 : romdata_int = 'h2822;
    'hc85 : romdata_int = 'h406e;
    'hc86 : romdata_int = 'h6e00;
    'hc87 : romdata_int = 'hd4b8;
    'hc88 : romdata_int = 'he600;
    'hc89 : romdata_int = 'hec5e;
    'hc8a : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc8b : romdata_int = 'h4f2;
    'hc8c : romdata_int = 'h120b;
    'hc8d : romdata_int = 'h5d0b;
    'hc8e : romdata_int = 'h7000;
    'hc8f : romdata_int = 'h7656;
    'hc90 : romdata_int = 'hc846;
    'hc91 : romdata_int = 'hda3a;
    'hc92 : romdata_int = 'he800;
    'hc93 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc94 : romdata_int = 'h701;
    'hc95 : romdata_int = 'h1447;
    'hc96 : romdata_int = 'h56b7;
    'hc97 : romdata_int = 'h6256;
    'hc98 : romdata_int = 'h7200;
    'hc99 : romdata_int = 'h7edf;
    'hc9a : romdata_int = 'ha6a7;
    'hc9b : romdata_int = 'hea00;
    'hc9c : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc9d : romdata_int = 'h832;
    'hc9e : romdata_int = 'haa2;
    'hc9f : romdata_int = 'h114b;
    'hca0 : romdata_int = 'h6840;
    'hca1 : romdata_int = 'h7400;
    'hca2 : romdata_int = 'h869c;
    'hca3 : romdata_int = 'hb229;
    'hca4 : romdata_int = 'hec00;
    'hca5 : romdata_int = 'h673c; // Line descriptor for 2_3
    'hca6 : romdata_int = 'h328;
    'hca7 : romdata_int = 'h648;
    'hca8 : romdata_int = 'h80a;
    'hca9 : romdata_int = 'h10f5;
    'hcaa : romdata_int = 'h7600;
    'hcab : romdata_int = 'hcb1e;
    'hcac : romdata_int = 'hdc17;
    'hcad : romdata_int = 'hee00;
    'hcae : romdata_int = 'hb2d; // Line descriptor for 3_4
    'hcaf : romdata_int = 'h0;
    'hcb0 : romdata_int = 'h534;
    'hcb1 : romdata_int = 'h69b;
    'hcb2 : romdata_int = 'hcd7;
    'hcb3 : romdata_int = 'h14c4;
    'hcb4 : romdata_int = 'h3e61;
    'hcb5 : romdata_int = 'h5a00;
    'hcb6 : romdata_int = 'h76bb;
    'hcb7 : romdata_int = 'h8a3b;
    'hcb8 : romdata_int = 'hb400;
    'hcb9 : romdata_int = 'hbcad;
    'hcba : romdata_int = 'hfd1a;
    'hcbb : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hcbc : romdata_int = 'h200;
    'hcbd : romdata_int = 'h651;
    'hcbe : romdata_int = 'he09;
    'hcbf : romdata_int = 'h122e;
    'hcc0 : romdata_int = 'h4f3e;
    'hcc1 : romdata_int = 'h50b5;
    'hcc2 : romdata_int = 'h5c00;
    'hcc3 : romdata_int = 'h7d0c;
    'hcc4 : romdata_int = 'ha4d1;
    'hcc5 : romdata_int = 'hb600;
    'hcc6 : romdata_int = 'he34b;
    'hcc7 : romdata_int = 'h102b4;
    'hcc8 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hcc9 : romdata_int = 'h296;
    'hcca : romdata_int = 'h400;
    'hccb : romdata_int = 'h50f;
    'hccc : romdata_int = 'hf52;
    'hccd : romdata_int = 'h3c46;
    'hcce : romdata_int = 'h515b;
    'hccf : romdata_int = 'h5e00;
    'hcd0 : romdata_int = 'h66b0;
    'hcd1 : romdata_int = 'hab47;
    'hcd2 : romdata_int = 'hb49d;
    'hcd3 : romdata_int = 'hb800;
    'hcd4 : romdata_int = 'he54c;
    'hcd5 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hcd6 : romdata_int = 'h600;
    'hcd7 : romdata_int = 'ha8c;
    'hcd8 : romdata_int = 'he58;
    'hcd9 : romdata_int = 'h100c;
    'hcda : romdata_int = 'h1135;
    'hcdb : romdata_int = 'h2323;
    'hcdc : romdata_int = 'h6000;
    'hcdd : romdata_int = 'h6106;
    'hcde : romdata_int = 'h649b;
    'hcdf : romdata_int = 'hba00;
    'hce0 : romdata_int = 'hf6a5;
    'hce1 : romdata_int = 'h10c40;
    'hce2 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hce3 : romdata_int = 'h541;
    'hce4 : romdata_int = 'h800;
    'hce5 : romdata_int = 'h149d;
    'hce6 : romdata_int = 'h175b;
    'hce7 : romdata_int = 'h3abf;
    'hce8 : romdata_int = 'h4829;
    'hce9 : romdata_int = 'h5a1c;
    'hcea : romdata_int = 'h5d18;
    'hceb : romdata_int = 'h6200;
    'hcec : romdata_int = 'hbc00;
    'hced : romdata_int = 'hc814;
    'hcee : romdata_int = 'hd6bd;
    'hcef : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hcf0 : romdata_int = 'ha1f;
    'hcf1 : romdata_int = 'ha00;
    'hcf2 : romdata_int = 'hb16;
    'hcf3 : romdata_int = 'h12a1;
    'hcf4 : romdata_int = 'h3c4d;
    'hcf5 : romdata_int = 'h4131;
    'hcf6 : romdata_int = 'h6400;
    'hcf7 : romdata_int = 'h9364;
    'hcf8 : romdata_int = 'h9b0d;
    'hcf9 : romdata_int = 'hbc1f;
    'hcfa : romdata_int = 'hbe00;
    'hcfb : romdata_int = 'h10750;
    'hcfc : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hcfd : romdata_int = 'hb3b;
    'hcfe : romdata_int = 'hc00;
    'hcff : romdata_int = 'h10cc;
    'hd00 : romdata_int = 'h120c;
    'hd01 : romdata_int = 'h18c2;
    'hd02 : romdata_int = 'h212a;
    'hd03 : romdata_int = 'h6046;
    'hd04 : romdata_int = 'h6600;
    'hd05 : romdata_int = 'hb28a;
    'hd06 : romdata_int = 'hc000;
    'hd07 : romdata_int = 'hc46b;
    'hd08 : romdata_int = 'hd43d;
    'hd09 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd0a : romdata_int = 'he00;
    'hd0b : romdata_int = 'h1319;
    'hd0c : romdata_int = 'h1a96;
    'hd0d : romdata_int = 'h1cb5;
    'hd0e : romdata_int = 'h26a0;
    'hd0f : romdata_int = 'h433b;
    'hd10 : romdata_int = 'h5e3c;
    'hd11 : romdata_int = 'h6800;
    'hd12 : romdata_int = 'h8457;
    'hd13 : romdata_int = 'hc200;
    'hd14 : romdata_int = 'hd8c6;
    'hd15 : romdata_int = 'hf72b;
    'hd16 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd17 : romdata_int = 'h824;
    'hd18 : romdata_int = 'h1000;
    'hd19 : romdata_int = 'h104f;
    'hd1a : romdata_int = 'h14e0;
    'hd1b : romdata_int = 'h1948;
    'hd1c : romdata_int = 'h2a62;
    'hd1d : romdata_int = 'h6a00;
    'hd1e : romdata_int = 'h6e27;
    'hd1f : romdata_int = 'hb2ab;
    'hd20 : romdata_int = 'hc0ab;
    'hd21 : romdata_int = 'hc400;
    'hd22 : romdata_int = 'he892;
    'hd23 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd24 : romdata_int = 'h333;
    'hd25 : romdata_int = 'h48e;
    'hd26 : romdata_int = 'h8f0;
    'hd27 : romdata_int = 'hc5a;
    'hd28 : romdata_int = 'h1200;
    'hd29 : romdata_int = 'h3b1d;
    'hd2a : romdata_int = 'h6c00;
    'hd2b : romdata_int = 'h720c;
    'hd2c : romdata_int = 'hae1a;
    'hd2d : romdata_int = 'hc600;
    'hd2e : romdata_int = 'hd90f;
    'hd2f : romdata_int = 'hde59;
    'hd30 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd31 : romdata_int = 'h354;
    'hd32 : romdata_int = 'h86c;
    'hd33 : romdata_int = 'h1293;
    'hd34 : romdata_int = 'h1400;
    'hd35 : romdata_int = 'h1851;
    'hd36 : romdata_int = 'h1a0b;
    'hd37 : romdata_int = 'h6e00;
    'hd38 : romdata_int = 'h7eb3;
    'hd39 : romdata_int = 'h9d58;
    'hd3a : romdata_int = 'hc709;
    'hd3b : romdata_int = 'hc800;
    'hd3c : romdata_int = 'hc828;
    'hd3d : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd3e : romdata_int = 'h12;
    'hd3f : romdata_int = 'ha78;
    'hd40 : romdata_int = 'h1080;
    'hd41 : romdata_int = 'h1600;
    'hd42 : romdata_int = 'h1f0a;
    'hd43 : romdata_int = 'h2ea8;
    'hd44 : romdata_int = 'h7000;
    'hd45 : romdata_int = 'h7026;
    'hd46 : romdata_int = 'h7314;
    'hd47 : romdata_int = 'hc239;
    'hd48 : romdata_int = 'hca00;
    'hd49 : romdata_int = 'hf510;
    'hd4a : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd4b : romdata_int = 'h48;
    'hd4c : romdata_int = 'h4b1;
    'hd4d : romdata_int = 'h1800;
    'hd4e : romdata_int = 'h186d;
    'hd4f : romdata_int = 'h1a3a;
    'hd50 : romdata_int = 'h3f35;
    'hd51 : romdata_int = 'h694f;
    'hd52 : romdata_int = 'h7200;
    'hd53 : romdata_int = 'h98d5;
    'hd54 : romdata_int = 'hb44d;
    'hd55 : romdata_int = 'hcc00;
    'hd56 : romdata_int = 'hd0ae;
    'hd57 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd58 : romdata_int = 'h8ce;
    'hd59 : romdata_int = 'h14cd;
    'hd5a : romdata_int = 'h162a;
    'hd5b : romdata_int = 'h1a00;
    'hd5c : romdata_int = 'h1ac6;
    'hd5d : romdata_int = 'h52f9;
    'hd5e : romdata_int = 'h6a70;
    'hd5f : romdata_int = 'h7400;
    'hd60 : romdata_int = 'h8827;
    'hd61 : romdata_int = 'hce00;
    'hd62 : romdata_int = 'hd667;
    'hd63 : romdata_int = 'hdd18;
    'hd64 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd65 : romdata_int = 'h706;
    'hd66 : romdata_int = 'h8d7;
    'hd67 : romdata_int = 'h1962;
    'hd68 : romdata_int = 'h1b26;
    'hd69 : romdata_int = 'h1c00;
    'hd6a : romdata_int = 'h2c3b;
    'hd6b : romdata_int = 'h6765;
    'hd6c : romdata_int = 'h7600;
    'hd6d : romdata_int = 'h7c1f;
    'hd6e : romdata_int = 'hd000;
    'hd6f : romdata_int = 'hd287;
    'hd70 : romdata_int = 'he8be;
    'hd71 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd72 : romdata_int = 'h81b;
    'hd73 : romdata_int = 'hf0b;
    'hd74 : romdata_int = 'h1492;
    'hd75 : romdata_int = 'h1e00;
    'hd76 : romdata_int = 'h2541;
    'hd77 : romdata_int = 'h3488;
    'hd78 : romdata_int = 'h7800;
    'hd79 : romdata_int = 'h8882;
    'hd7a : romdata_int = 'had55;
    'hd7b : romdata_int = 'hcc4f;
    'hd7c : romdata_int = 'hd200;
    'hd7d : romdata_int = 'hfa38;
    'hd7e : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd7f : romdata_int = 'h6a2;
    'hd80 : romdata_int = 'hc67;
    'hd81 : romdata_int = 'hcc4;
    'hd82 : romdata_int = 'h12d9;
    'hd83 : romdata_int = 'h2000;
    'hd84 : romdata_int = 'h4675;
    'hd85 : romdata_int = 'h7a00;
    'hd86 : romdata_int = 'ha8bd;
    'hd87 : romdata_int = 'haabc;
    'hd88 : romdata_int = 'hb657;
    'hd89 : romdata_int = 'hd400;
    'hd8a : romdata_int = 'he49e;
    'hd8b : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd8c : romdata_int = 'h550;
    'hd8d : romdata_int = 'h727;
    'hd8e : romdata_int = 'h73e;
    'hd8f : romdata_int = 'h2200;
    'hd90 : romdata_int = 'h38c0;
    'hd91 : romdata_int = 'h4eaa;
    'hd92 : romdata_int = 'h7c00;
    'hd93 : romdata_int = 'h8b4c;
    'hd94 : romdata_int = 'hb034;
    'hd95 : romdata_int = 'hccfb;
    'hd96 : romdata_int = 'hd600;
    'hd97 : romdata_int = 'h102e2;
    'hd98 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd99 : romdata_int = 'hce4;
    'hd9a : romdata_int = 'hce6;
    'hd9b : romdata_int = 'hecb;
    'hd9c : romdata_int = 'h16f0;
    'hd9d : romdata_int = 'h1d41;
    'hd9e : romdata_int = 'h2400;
    'hd9f : romdata_int = 'h6538;
    'hda0 : romdata_int = 'h78d9;
    'hda1 : romdata_int = 'h7e00;
    'hda2 : romdata_int = 'hd800;
    'hda3 : romdata_int = 'hef34;
    'hda4 : romdata_int = 'hf2ff;
    'hda5 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hda6 : romdata_int = 'h2fc;
    'hda7 : romdata_int = 'h944;
    'hda8 : romdata_int = 'h182f;
    'hda9 : romdata_int = 'h1b5a;
    'hdaa : romdata_int = 'h2600;
    'hdab : romdata_int = 'h474e;
    'hdac : romdata_int = 'h8000;
    'hdad : romdata_int = 'h9b56;
    'hdae : romdata_int = 'haeb0;
    'hdaf : romdata_int = 'hc037;
    'hdb0 : romdata_int = 'hda00;
    'hdb1 : romdata_int = 'hfecf;
    'hdb2 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hdb3 : romdata_int = 'hb35;
    'hdb4 : romdata_int = 'h1013;
    'hdb5 : romdata_int = 'h14f6;
    'hdb6 : romdata_int = 'h2800;
    'hdb7 : romdata_int = 'h36a6;
    'hdb8 : romdata_int = 'h4c87;
    'hdb9 : romdata_int = 'h5cdd;
    'hdba : romdata_int = 'h8200;
    'hdbb : romdata_int = 'h9467;
    'hdbc : romdata_int = 'hdc00;
    'hdbd : romdata_int = 'he226;
    'hdbe : romdata_int = 'h10941;
    'hdbf : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hdc0 : romdata_int = 'h22c;
    'hdc1 : romdata_int = 'h48c;
    'hdc2 : romdata_int = 'h8a9;
    'hdc3 : romdata_int = 'h16f5;
    'hdc4 : romdata_int = 'h2099;
    'hdc5 : romdata_int = 'h2a00;
    'hdc6 : romdata_int = 'h70b4;
    'hdc7 : romdata_int = 'h8400;
    'hdc8 : romdata_int = 'ha46a;
    'hdc9 : romdata_int = 'hcf4b;
    'hdca : romdata_int = 'hdc62;
    'hdcb : romdata_int = 'hde00;
    'hdcc : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hdcd : romdata_int = 'h3c;
    'hdce : romdata_int = 'h52e;
    'hdcf : romdata_int = 'h8fd;
    'hdd0 : romdata_int = 'h1085;
    'hdd1 : romdata_int = 'h12a2;
    'hdd2 : romdata_int = 'h2c00;
    'hdd3 : romdata_int = 'h8600;
    'hdd4 : romdata_int = 'ha2b7;
    'hdd5 : romdata_int = 'ha83e;
    'hdd6 : romdata_int = 'hc55c;
    'hdd7 : romdata_int = 'he000;
    'hdd8 : romdata_int = 'hf107;
    'hdd9 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hdda : romdata_int = 'h74;
    'hddb : romdata_int = 'haa3;
    'hddc : romdata_int = 'hcae;
    'hddd : romdata_int = 'h2e00;
    'hdde : romdata_int = 'h2ec8;
    'hddf : romdata_int = 'h4818;
    'hde0 : romdata_int = 'h6f57;
    'hde1 : romdata_int = 'h80bb;
    'hde2 : romdata_int = 'h8800;
    'hde3 : romdata_int = 'hd457;
    'hde4 : romdata_int = 'hdb14;
    'hde5 : romdata_int = 'he200;
    'hde6 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hde7 : romdata_int = 'h129;
    'hde8 : romdata_int = 'h124b;
    'hde9 : romdata_int = 'h1748;
    'hdea : romdata_int = 'h3000;
    'hdeb : romdata_int = 'h3743;
    'hdec : romdata_int = 'h4cd6;
    'hded : romdata_int = 'h8a00;
    'hdee : romdata_int = 'h9cc2;
    'hdef : romdata_int = 'ha159;
    'hdf0 : romdata_int = 'he400;
    'hdf1 : romdata_int = 'hf923;
    'hdf2 : romdata_int = 'h10af7;
    'hdf3 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hdf4 : romdata_int = 'h108a;
    'hdf5 : romdata_int = 'h126a;
    'hdf6 : romdata_int = 'h1700;
    'hdf7 : romdata_int = 'h2d36;
    'hdf8 : romdata_int = 'h3200;
    'hdf9 : romdata_int = 'h552f;
    'hdfa : romdata_int = 'h8c00;
    'hdfb : romdata_int = 'h9f54;
    'hdfc : romdata_int = 'ha242;
    'hdfd : romdata_int = 'hb8aa;
    'hdfe : romdata_int = 'he600;
    'hdff : romdata_int = 'hed1c;
    'he00 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he01 : romdata_int = 'haf;
    'he02 : romdata_int = 'hf0f;
    'he03 : romdata_int = 'h1c43;
    'he04 : romdata_int = 'h1c91;
    'he05 : romdata_int = 'h32a1;
    'he06 : romdata_int = 'h3400;
    'he07 : romdata_int = 'h749d;
    'he08 : romdata_int = 'h8655;
    'he09 : romdata_int = 'h8e00;
    'he0a : romdata_int = 'he800;
    'he0b : romdata_int = 'hf0f8;
    'he0c : romdata_int = 'h10155;
    'he0d : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he0e : romdata_int = 'hcb1;
    'he0f : romdata_int = 'h113b;
    'he10 : romdata_int = 'h126d;
    'he11 : romdata_int = 'h2849;
    'he12 : romdata_int = 'h3600;
    'he13 : romdata_int = 'h4524;
    'he14 : romdata_int = 'h5eb6;
    'he15 : romdata_int = 'h9000;
    'he16 : romdata_int = 'h92a9;
    'he17 : romdata_int = 'hc2af;
    'he18 : romdata_int = 'hea00;
    'he19 : romdata_int = 'hec06;
    'he1a : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he1b : romdata_int = 'h149f;
    'he1c : romdata_int = 'h1cc2;
    'he1d : romdata_int = 'h1d5d;
    'he1e : romdata_int = 'h329e;
    'he1f : romdata_int = 'h3800;
    'he20 : romdata_int = 'h56be;
    'he21 : romdata_int = 'h8e5f;
    'he22 : romdata_int = 'h9200;
    'he23 : romdata_int = 'h9723;
    'he24 : romdata_int = 'he0bc;
    'he25 : romdata_int = 'hec00;
    'he26 : romdata_int = 'h10137;
    'he27 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he28 : romdata_int = 'h37;
    'he29 : romdata_int = 'ha7e;
    'he2a : romdata_int = 'h1602;
    'he2b : romdata_int = 'h1820;
    'he2c : romdata_int = 'h242c;
    'he2d : romdata_int = 'h3a00;
    'he2e : romdata_int = 'h6221;
    'he2f : romdata_int = 'h9400;
    'he30 : romdata_int = 'ha040;
    'he31 : romdata_int = 'hb91e;
    'he32 : romdata_int = 'hd0aa;
    'he33 : romdata_int = 'hee00;
    'he34 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he35 : romdata_int = 'h622;
    'he36 : romdata_int = 'hc4b;
    'he37 : romdata_int = 'hc84;
    'he38 : romdata_int = 'h14a5;
    'he39 : romdata_int = 'h2857;
    'he3a : romdata_int = 'h3c00;
    'he3b : romdata_int = 'h8339;
    'he3c : romdata_int = 'h8c7b;
    'he3d : romdata_int = 'h9600;
    'he3e : romdata_int = 'hb733;
    'he3f : romdata_int = 'hf000;
    'he40 : romdata_int = 'hfc8f;
    'he41 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he42 : romdata_int = 'h144;
    'he43 : romdata_int = 'h952;
    'he44 : romdata_int = 'he62;
    'he45 : romdata_int = 'h1a5d;
    'he46 : romdata_int = 'h3e00;
    'he47 : romdata_int = 'h583b;
    'he48 : romdata_int = 'h761f;
    'he49 : romdata_int = 'h8f18;
    'he4a : romdata_int = 'h9800;
    'he4b : romdata_int = 'hc6e7;
    'he4c : romdata_int = 'hf200;
    'he4d : romdata_int = 'h10d42;
    'he4e : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he4f : romdata_int = 'h2fd;
    'he50 : romdata_int = 'h4ae;
    'he51 : romdata_int = 'h654;
    'he52 : romdata_int = 'h104d;
    'he53 : romdata_int = 'h2328;
    'he54 : romdata_int = 'h4000;
    'he55 : romdata_int = 'h5a16;
    'he56 : romdata_int = 'h8c8c;
    'he57 : romdata_int = 'h9a00;
    'he58 : romdata_int = 'hee94;
    'he59 : romdata_int = 'hf400;
    'he5a : romdata_int = 'hfe98;
    'he5b : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he5c : romdata_int = 'h14e1;
    'he5d : romdata_int = 'h1cf8;
    'he5e : romdata_int = 'h1d4f;
    'he5f : romdata_int = 'h4200;
    'he60 : romdata_int = 'h4a2d;
    'he61 : romdata_int = 'h548a;
    'he62 : romdata_int = 'h690d;
    'he63 : romdata_int = 'h821c;
    'he64 : romdata_int = 'h9c00;
    'he65 : romdata_int = 'hbecc;
    'he66 : romdata_int = 'hf600;
    'he67 : romdata_int = 'h1046b;
    'he68 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he69 : romdata_int = 'h52a;
    'he6a : romdata_int = 'hea5;
    'he6b : romdata_int = 'h1960;
    'he6c : romdata_int = 'h4400;
    'he6d : romdata_int = 'h4436;
    'he6e : romdata_int = 'h4a17;
    'he6f : romdata_int = 'h745b;
    'he70 : romdata_int = 'h7afb;
    'he71 : romdata_int = 'h9e00;
    'he72 : romdata_int = 'hd322;
    'he73 : romdata_int = 'hda7f;
    'he74 : romdata_int = 'hf800;
    'he75 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he76 : romdata_int = 'h680;
    'he77 : romdata_int = 'ha23;
    'he78 : romdata_int = 'h1604;
    'he79 : romdata_int = 'h1d1d;
    'he7a : romdata_int = 'h352f;
    'he7b : romdata_int = 'h4600;
    'he7c : romdata_int = 'h6a8f;
    'he7d : romdata_int = 'ha000;
    'he7e : romdata_int = 'hacad;
    'he7f : romdata_int = 'he133;
    'he80 : romdata_int = 'hf566;
    'he81 : romdata_int = 'hfa00;
    'he82 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he83 : romdata_int = 'h6ae;
    'he84 : romdata_int = 'hb60;
    'he85 : romdata_int = 'hd54;
    'he86 : romdata_int = 'h1ab8;
    'he87 : romdata_int = 'h3836;
    'he88 : romdata_int = 'h4800;
    'he89 : romdata_int = 'h8533;
    'he8a : romdata_int = 'h9ea4;
    'he8b : romdata_int = 'ha200;
    'he8c : romdata_int = 'hea08;
    'he8d : romdata_int = 'hf942;
    'he8e : romdata_int = 'hfc00;
    'he8f : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he90 : romdata_int = 'h31b;
    'he91 : romdata_int = 'h1247;
    'he92 : romdata_int = 'h183b;
    'he93 : romdata_int = 'h1ab0;
    'he94 : romdata_int = 'h1c6b;
    'he95 : romdata_int = 'h4a00;
    'he96 : romdata_int = 'h6d4b;
    'he97 : romdata_int = 'h9936;
    'he98 : romdata_int = 'ha400;
    'he99 : romdata_int = 'hcafb;
    'he9a : romdata_int = 'hfe00;
    'he9b : romdata_int = 'h10a72;
    'he9c : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he9d : romdata_int = 'hf19;
    'he9e : romdata_int = 'h140a;
    'he9f : romdata_int = 'h1d2f;
    'hea0 : romdata_int = 'h2a8a;
    'hea1 : romdata_int = 'h42f3;
    'hea2 : romdata_int = 'h4c00;
    'hea3 : romdata_int = 'h8040;
    'hea4 : romdata_int = 'ha600;
    'hea5 : romdata_int = 'hb0c0;
    'hea6 : romdata_int = 'hfaf9;
    'hea7 : romdata_int = 'h10000;
    'hea8 : romdata_int = 'h10509;
    'hea9 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'heaa : romdata_int = 'ha3;
    'heab : romdata_int = 'he2e;
    'heac : romdata_int = 'h1523;
    'head : romdata_int = 'h265f;
    'heae : romdata_int = 'h4085;
    'heaf : romdata_int = 'h4e00;
    'heb0 : romdata_int = 'h6207;
    'heb1 : romdata_int = 'ha66b;
    'heb2 : romdata_int = 'ha800;
    'heb3 : romdata_int = 'hcacd;
    'heb4 : romdata_int = 'hde1d;
    'heb5 : romdata_int = 'h10200;
    'heb6 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'heb7 : romdata_int = 'h8d;
    'heb8 : romdata_int = 'hf8;
    'heb9 : romdata_int = 'h16eb;
    'heba : romdata_int = 'h189e;
    'hebb : romdata_int = 'h1a54;
    'hebc : romdata_int = 'h5000;
    'hebd : romdata_int = 'h7a8b;
    'hebe : romdata_int = 'h8658;
    'hebf : romdata_int = 'haa00;
    'hec0 : romdata_int = 'hce3a;
    'hec1 : romdata_int = 'hf33f;
    'hec2 : romdata_int = 'h10400;
    'hec3 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hec4 : romdata_int = 'had1;
    'hec5 : romdata_int = 'h10ba;
    'hec6 : romdata_int = 'h16b0;
    'hec7 : romdata_int = 'h1a11;
    'hec8 : romdata_int = 'h5200;
    'hec9 : romdata_int = 'h5904;
    'heca : romdata_int = 'h910f;
    'hecb : romdata_int = 'ha6f6;
    'hecc : romdata_int = 'hac00;
    'hecd : romdata_int = 'hbe82;
    'hece : romdata_int = 'h10600;
    'hecf : romdata_int = 'h108b2;
    'hed0 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hed1 : romdata_int = 'h207;
    'hed2 : romdata_int = 'h212;
    'hed3 : romdata_int = 'h6c2;
    'hed4 : romdata_int = 'h3041;
    'hed5 : romdata_int = 'h313a;
    'hed6 : romdata_int = 'h5400;
    'hed7 : romdata_int = 'h6d19;
    'hed8 : romdata_int = 'h7ec9;
    'hed9 : romdata_int = 'hae00;
    'heda : romdata_int = 'hbab5;
    'hedb : romdata_int = 'hea6d;
    'hedc : romdata_int = 'h10800;
    'hedd : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hede : romdata_int = 'h23b;
    'hedf : romdata_int = 'h425;
    'hee0 : romdata_int = 'h82e;
    'hee1 : romdata_int = 'h16a7;
    'hee2 : romdata_int = 'h5265;
    'hee3 : romdata_int = 'h5600;
    'hee4 : romdata_int = 'h9102;
    'hee5 : romdata_int = 'h9539;
    'hee6 : romdata_int = 'hb000;
    'hee7 : romdata_int = 'he6c4;
    'hee8 : romdata_int = 'he74c;
    'hee9 : romdata_int = 'h10a00;
    'heea : romdata_int = 'h6b2d; // Line descriptor for 3_4
    'heeb : romdata_int = 'h2a0;
    'heec : romdata_int = 'he0d;
    'heed : romdata_int = 'h1871;
    'heee : romdata_int = 'h1e45;
    'heef : romdata_int = 'h56ae;
    'hef0 : romdata_int = 'h5800;
    'hef1 : romdata_int = 'h78a8;
    'hef2 : romdata_int = 'h96d4;
    'hef3 : romdata_int = 'hb200;
    'hef4 : romdata_int = 'hba26;
    'hef5 : romdata_int = 'h10687;
    'hef6 : romdata_int = 'h10c00;
    'hef7 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hef8 : romdata_int = 'h0;
    'hef9 : romdata_int = 'hc68;
    'hefa : romdata_int = 'h1945;
    'hefb : romdata_int = 'h1eb5;
    'hefc : romdata_int = 'h1f3f;
    'hefd : romdata_int = 'h22f3;
    'hefe : romdata_int = 'h3279;
    'heff : romdata_int = 'h4800;
    'hf00 : romdata_int = 'h4e3d;
    'hf01 : romdata_int = 'h6248;
    'hf02 : romdata_int = 'h9000;
    'hf03 : romdata_int = 'ha222;
    'hf04 : romdata_int = 'hacc8;
    'hf05 : romdata_int = 'hd800;
    'hf06 : romdata_int = 'hfae7;
    'hf07 : romdata_int = 'h11702;
    'hf08 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf09 : romdata_int = 'h200;
    'hf0a : romdata_int = 'h1207;
    'hf0b : romdata_int = 'h14f2;
    'hf0c : romdata_int = 'h1c60;
    'hf0d : romdata_int = 'h233b;
    'hf0e : romdata_int = 'h374a;
    'hf0f : romdata_int = 'h4321;
    'hf10 : romdata_int = 'h4a00;
    'hf11 : romdata_int = 'h5329;
    'hf12 : romdata_int = 'h7e61;
    'hf13 : romdata_int = 'h9200;
    'hf14 : romdata_int = 'hc017;
    'hf15 : romdata_int = 'hc567;
    'hf16 : romdata_int = 'hda00;
    'hf17 : romdata_int = 'hed58;
    'hf18 : romdata_int = 'hf2d3;
    'hf19 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf1a : romdata_int = 'h400;
    'hf1b : romdata_int = 'ha5f;
    'hf1c : romdata_int = 'he1f;
    'hf1d : romdata_int = 'h14da;
    'hf1e : romdata_int = 'h186b;
    'hf1f : romdata_int = 'h261c;
    'hf20 : romdata_int = 'h2b55;
    'hf21 : romdata_int = 'h4c00;
    'hf22 : romdata_int = 'h614c;
    'hf23 : romdata_int = 'h863a;
    'hf24 : romdata_int = 'h9400;
    'hf25 : romdata_int = 'h9c9c;
    'hf26 : romdata_int = 'hd4e2;
    'hf27 : romdata_int = 'hdc00;
    'hf28 : romdata_int = 'hed4d;
    'hf29 : romdata_int = 'hfab7;
    'hf2a : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf2b : romdata_int = 'h600;
    'hf2c : romdata_int = 'ha1c;
    'hf2d : romdata_int = 'ha3b;
    'hf2e : romdata_int = 'h1241;
    'hf2f : romdata_int = 'h16fe;
    'hf30 : romdata_int = 'h1e4c;
    'hf31 : romdata_int = 'h251a;
    'hf32 : romdata_int = 'h4e00;
    'hf33 : romdata_int = 'h50d1;
    'hf34 : romdata_int = 'h74d8;
    'hf35 : romdata_int = 'h9089;
    'hf36 : romdata_int = 'h9600;
    'hf37 : romdata_int = 'hbcb8;
    'hf38 : romdata_int = 'hde00;
    'hf39 : romdata_int = 'h10007;
    'hf3a : romdata_int = 'h102a2;
    'hf3b : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf3c : romdata_int = 'h800;
    'hf3d : romdata_int = 'h94d;
    'hf3e : romdata_int = 'hc1a;
    'hf3f : romdata_int = 'heb4;
    'hf40 : romdata_int = 'h1eb8;
    'hf41 : romdata_int = 'h3c3e;
    'hf42 : romdata_int = 'h3eb0;
    'hf43 : romdata_int = 'h5000;
    'hf44 : romdata_int = 'h62ce;
    'hf45 : romdata_int = 'h6ca7;
    'hf46 : romdata_int = 'h9800;
    'hf47 : romdata_int = 'ha85a;
    'hf48 : romdata_int = 'hd011;
    'hf49 : romdata_int = 'he000;
    'hf4a : romdata_int = 'hf403;
    'hf4b : romdata_int = 'h10d0e;
    'hf4c : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf4d : romdata_int = 'h4;
    'hf4e : romdata_int = 'ha00;
    'hf4f : romdata_int = 'ha71;
    'hf50 : romdata_int = 'h127d;
    'hf51 : romdata_int = 'h1b3e;
    'hf52 : romdata_int = 'h20e5;
    'hf53 : romdata_int = 'h2c7a;
    'hf54 : romdata_int = 'h5200;
    'hf55 : romdata_int = 'h58df;
    'hf56 : romdata_int = 'h6613;
    'hf57 : romdata_int = 'h9a00;
    'hf58 : romdata_int = 'hc23d;
    'hf59 : romdata_int = 'hd30f;
    'hf5a : romdata_int = 'he200;
    'hf5b : romdata_int = 'h10003;
    'hf5c : romdata_int = 'h102ac;
    'hf5d : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf5e : romdata_int = 'hc00;
    'hf5f : romdata_int = 'heda;
    'hf60 : romdata_int = 'h10ea;
    'hf61 : romdata_int = 'h163f;
    'hf62 : romdata_int = 'h16a8;
    'hf63 : romdata_int = 'h1a45;
    'hf64 : romdata_int = 'h3646;
    'hf65 : romdata_int = 'h5400;
    'hf66 : romdata_int = 'h544b;
    'hf67 : romdata_int = 'h726f;
    'hf68 : romdata_int = 'h9c00;
    'hf69 : romdata_int = 'hb03d;
    'hf6a : romdata_int = 'hb156;
    'hf6b : romdata_int = 'he400;
    'hf6c : romdata_int = 'h10898;
    'hf6d : romdata_int = 'h10f40;
    'hf6e : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf6f : romdata_int = 'h94f;
    'hf70 : romdata_int = 'hc4e;
    'hf71 : romdata_int = 'he00;
    'hf72 : romdata_int = 'h14bc;
    'hf73 : romdata_int = 'h14e3;
    'hf74 : romdata_int = 'h1caf;
    'hf75 : romdata_int = 'h2723;
    'hf76 : romdata_int = 'h5600;
    'hf77 : romdata_int = 'h5a7b;
    'hf78 : romdata_int = 'h7e44;
    'hf79 : romdata_int = 'h9275;
    'hf7a : romdata_int = 'h9e00;
    'hf7b : romdata_int = 'hac5b;
    'hf7c : romdata_int = 'he600;
    'hf7d : romdata_int = 'he8ce;
    'hf7e : romdata_int = 'h11108;
    'hf7f : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf80 : romdata_int = 'he1;
    'hf81 : romdata_int = 'h1000;
    'hf82 : romdata_int = 'h1106;
    'hf83 : romdata_int = 'h122b;
    'hf84 : romdata_int = 'h14f8;
    'hf85 : romdata_int = 'h1c69;
    'hf86 : romdata_int = 'h28f7;
    'hf87 : romdata_int = 'h5800;
    'hf88 : romdata_int = 'h6824;
    'hf89 : romdata_int = 'h8cec;
    'hf8a : romdata_int = 'h9af9;
    'hf8b : romdata_int = 'ha000;
    'hf8c : romdata_int = 'hc8a5;
    'hf8d : romdata_int = 'he060;
    'hf8e : romdata_int = 'he800;
    'hf8f : romdata_int = 'h10a3b;
    'hf90 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf91 : romdata_int = 'hec;
    'hf92 : romdata_int = 'h31e;
    'hf93 : romdata_int = 'h49a;
    'hf94 : romdata_int = 'h523;
    'hf95 : romdata_int = 'h1200;
    'hf96 : romdata_int = 'h1aa2;
    'hf97 : romdata_int = 'h34c6;
    'hf98 : romdata_int = 'h490b;
    'hf99 : romdata_int = 'h5a00;
    'hf9a : romdata_int = 'h786e;
    'hf9b : romdata_int = 'ha200;
    'hf9c : romdata_int = 'hc6f3;
    'hf9d : romdata_int = 'hd520;
    'hf9e : romdata_int = 'hea00;
    'hf9f : romdata_int = 'hf6dd;
    'hfa0 : romdata_int = 'h11e9a;
    'hfa1 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hfa2 : romdata_int = 'h65a;
    'hfa3 : romdata_int = 'h8ab;
    'hfa4 : romdata_int = 'h1400;
    'hfa5 : romdata_int = 'h183c;
    'hfa6 : romdata_int = 'h186e;
    'hfa7 : romdata_int = 'h1b4c;
    'hfa8 : romdata_int = 'h3308;
    'hfa9 : romdata_int = 'h5c00;
    'hfaa : romdata_int = 'h5eb6;
    'hfab : romdata_int = 'h82b7;
    'hfac : romdata_int = 'ha2f6;
    'hfad : romdata_int = 'ha400;
    'hfae : romdata_int = 'hb91e;
    'hfaf : romdata_int = 'hec00;
    'hfb0 : romdata_int = 'hf11a;
    'hfb1 : romdata_int = 'hf428;
    'hfb2 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hfb3 : romdata_int = 'h1072;
    'hfb4 : romdata_int = 'h10ee;
    'hfb5 : romdata_int = 'h1600;
    'hfb6 : romdata_int = 'h1966;
    'hfb7 : romdata_int = 'h1e0f;
    'hfb8 : romdata_int = 'h1f50;
    'hfb9 : romdata_int = 'h4344;
    'hfba : romdata_int = 'h5e00;
    'hfbb : romdata_int = 'h707b;
    'hfbc : romdata_int = 'h833f;
    'hfbd : romdata_int = 'h9697;
    'hfbe : romdata_int = 'ha600;
    'hfbf : romdata_int = 'hb50a;
    'hfc0 : romdata_int = 'hee00;
    'hfc1 : romdata_int = 'hfcfa;
    'hfc2 : romdata_int = 'h11156;
    'hfc3 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hfc4 : romdata_int = 'hb;
    'hfc5 : romdata_int = 'h164;
    'hfc6 : romdata_int = 'h44e;
    'hfc7 : romdata_int = 'h142f;
    'hfc8 : romdata_int = 'h16f5;
    'hfc9 : romdata_int = 'h1800;
    'hfca : romdata_int = 'h3cf2;
    'hfcb : romdata_int = 'h5d00;
    'hfcc : romdata_int = 'h6000;
    'hfcd : romdata_int = 'h7a79;
    'hfce : romdata_int = 'ha0f6;
    'hfcf : romdata_int = 'ha800;
    'hfd0 : romdata_int = 'haaa2;
    'hfd1 : romdata_int = 'he2c1;
    'hfd2 : romdata_int = 'hf000;
    'hfd3 : romdata_int = 'h10c26;
    'hfd4 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hfd5 : romdata_int = 'h60e;
    'hfd6 : romdata_int = 'h88f;
    'hfd7 : romdata_int = 'he7e;
    'hfd8 : romdata_int = 'h129d;
    'hfd9 : romdata_int = 'h1a00;
    'hfda : romdata_int = 'h2032;
    'hfdb : romdata_int = 'h3b2f;
    'hfdc : romdata_int = 'h6200;
    'hfdd : romdata_int = 'h870b;
    'hfde : romdata_int = 'h8c33;
    'hfdf : romdata_int = 'h9859;
    'hfe0 : romdata_int = 'ha67a;
    'hfe1 : romdata_int = 'haa00;
    'hfe2 : romdata_int = 'hd8ca;
    'hfe3 : romdata_int = 'hf200;
    'hfe4 : romdata_int = 'h10661;
    'hfe5 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hfe6 : romdata_int = 'he23;
    'hfe7 : romdata_int = 'h174b;
    'hfe8 : romdata_int = 'h1c00;
    'hfe9 : romdata_int = 'h1ee2;
    'hfea : romdata_int = 'h223a;
    'hfeb : romdata_int = 'h2cc4;
    'hfec : romdata_int = 'h40ee;
    'hfed : romdata_int = 'h6400;
    'hfee : romdata_int = 'h7c94;
    'hfef : romdata_int = 'h8a63;
    'hff0 : romdata_int = 'ha607;
    'hff1 : romdata_int = 'hac00;
    'hff2 : romdata_int = 'haf39;
    'hff3 : romdata_int = 'hf400;
    'hff4 : romdata_int = 'hff05;
    'hff5 : romdata_int = 'h10566;
    'hff6 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hff7 : romdata_int = 'h683;
    'hff8 : romdata_int = 'hac5;
    'hff9 : romdata_int = 'he70;
    'hffa : romdata_int = 'hf46;
    'hffb : romdata_int = 'h16fc;
    'hffc : romdata_int = 'h18cb;
    'hffd : romdata_int = 'h1e00;
    'hffe : romdata_int = 'h6600;
    'hfff : romdata_int = 'h7309;
    'h1000: romdata_int = 'h8883;
    'h1001: romdata_int = 'hae00;
    'h1002: romdata_int = 'hc63b;
    'h1003: romdata_int = 'hd6a1;
    'h1004: romdata_int = 'hdee7;
    'h1005: romdata_int = 'hf225;
    'h1006: romdata_int = 'hf600;
    'h1007: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h1008: romdata_int = 'h137;
    'h1009: romdata_int = 'ha67;
    'h100a: romdata_int = 'hd2c;
    'h100b: romdata_int = 'h1745;
    'h100c: romdata_int = 'h1e47;
    'h100d: romdata_int = 'h2000;
    'h100e: romdata_int = 'h22ba;
    'h100f: romdata_int = 'h6800;
    'h1010: romdata_int = 'h7caf;
    'h1011: romdata_int = 'h8a48;
    'h1012: romdata_int = 'h9d5a;
    'h1013: romdata_int = 'hb000;
    'h1014: romdata_int = 'hc94d;
    'h1015: romdata_int = 'hf800;
    'h1016: romdata_int = 'h11a07;
    'h1017: romdata_int = 'h11ec5;
    'h1018: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h1019: romdata_int = 'h26b;
    'h101a: romdata_int = 'h261;
    'h101b: romdata_int = 'h291;
    'h101c: romdata_int = 'hd41;
    'h101d: romdata_int = 'h100b;
    'h101e: romdata_int = 'h2200;
    'h101f: romdata_int = 'h2298;
    'h1020: romdata_int = 'h5c73;
    'h1021: romdata_int = 'h6a00;
    'h1022: romdata_int = 'h8840;
    'h1023: romdata_int = 'h9e28;
    'h1024: romdata_int = 'hb200;
    'h1025: romdata_int = 'hc10d;
    'h1026: romdata_int = 'hf8cd;
    'h1027: romdata_int = 'hf8f8;
    'h1028: romdata_int = 'hfa00;
    'h1029: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h102a: romdata_int = 'h116;
    'h102b: romdata_int = 'h1158;
    'h102c: romdata_int = 'h12fd;
    'h102d: romdata_int = 'h18e5;
    'h102e: romdata_int = 'h20b5;
    'h102f: romdata_int = 'h2400;
    'h1030: romdata_int = 'h4658;
    'h1031: romdata_int = 'h6b4b;
    'h1032: romdata_int = 'h6c00;
    'h1033: romdata_int = 'h7629;
    'h1034: romdata_int = 'hb400;
    'h1035: romdata_int = 'hbb33;
    'h1036: romdata_int = 'hd0c6;
    'h1037: romdata_int = 'hf6eb;
    'h1038: romdata_int = 'hfc00;
    'h1039: romdata_int = 'hfeab;
    'h103a: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h103b: romdata_int = 'h4d8;
    'h103c: romdata_int = 'h825;
    'h103d: romdata_int = 'ha9f;
    'h103e: romdata_int = 'h1697;
    'h103f: romdata_int = 'h2080;
    'h1040: romdata_int = 'h2600;
    'h1041: romdata_int = 'h2b1c;
    'h1042: romdata_int = 'h4c87;
    'h1043: romdata_int = 'h6d09;
    'h1044: romdata_int = 'h6e00;
    'h1045: romdata_int = 'ha4e8;
    'h1046: romdata_int = 'hb600;
    'h1047: romdata_int = 'hc232;
    'h1048: romdata_int = 'hdcfa;
    'h1049: romdata_int = 'hef0e;
    'h104a: romdata_int = 'hfe00;
    'h104b: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h104c: romdata_int = 'h452;
    'h104d: romdata_int = 'h550;
    'h104e: romdata_int = 'h677;
    'h104f: romdata_int = 'h1cdd;
    'h1050: romdata_int = 'h2251;
    'h1051: romdata_int = 'h2800;
    'h1052: romdata_int = 'h3a54;
    'h1053: romdata_int = 'h4e09;
    'h1054: romdata_int = 'h6819;
    'h1055: romdata_int = 'h7000;
    'h1056: romdata_int = 'h9e23;
    'h1057: romdata_int = 'hb800;
    'h1058: romdata_int = 'hd6d3;
    'h1059: romdata_int = 'heae1;
    'h105a: romdata_int = 'h10000;
    'h105b: romdata_int = 'h11655;
    'h105c: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h105d: romdata_int = 'h328;
    'h105e: romdata_int = 'h1b37;
    'h105f: romdata_int = 'h1ca6;
    'h1060: romdata_int = 'h1cd6;
    'h1061: romdata_int = 'h2359;
    'h1062: romdata_int = 'h2a00;
    'h1063: romdata_int = 'h351d;
    'h1064: romdata_int = 'h7074;
    'h1065: romdata_int = 'h7200;
    'h1066: romdata_int = 'h792a;
    'h1067: romdata_int = 'h9a12;
    'h1068: romdata_int = 'hb94e;
    'h1069: romdata_int = 'hba00;
    'h106a: romdata_int = 'he89b;
    'h106b: romdata_int = 'h10200;
    'h106c: romdata_int = 'h10679;
    'h106d: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h106e: romdata_int = 'h20d;
    'h106f: romdata_int = 'hd08;
    'h1070: romdata_int = 'hd3f;
    'h1071: romdata_int = 'h20a8;
    'h1072: romdata_int = 'h2067;
    'h1073: romdata_int = 'h2149;
    'h1074: romdata_int = 'h2c00;
    'h1075: romdata_int = 'h56a6;
    'h1076: romdata_int = 'h5a86;
    'h1077: romdata_int = 'h7400;
    'h1078: romdata_int = 'h96c1;
    'h1079: romdata_int = 'h989c;
    'h107a: romdata_int = 'hbc00;
    'h107b: romdata_int = 'hde7a;
    'h107c: romdata_int = 'h10400;
    'h107d: romdata_int = 'h114fa;
    'h107e: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h107f: romdata_int = 'h841;
    'h1080: romdata_int = 'h952;
    'h1081: romdata_int = 'hf3f;
    'h1082: romdata_int = 'he90;
    'h1083: romdata_int = 'hf63;
    'h1084: romdata_int = 'h2e00;
    'h1085: romdata_int = 'h44b3;
    'h1086: romdata_int = 'h54bb;
    'h1087: romdata_int = 'h7600;
    'h1088: romdata_int = 'h7a60;
    'h1089: romdata_int = 'hb27d;
    'h108a: romdata_int = 'hbe00;
    'h108b: romdata_int = 'hca58;
    'h108c: romdata_int = 'he238;
    'h108d: romdata_int = 'h10600;
    'h108e: romdata_int = 'h112e4;
    'h108f: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h1090: romdata_int = 'hb0;
    'h1091: romdata_int = 'h40f;
    'h1092: romdata_int = 'habd;
    'h1093: romdata_int = 'hb32;
    'h1094: romdata_int = 'h1678;
    'h1095: romdata_int = 'h1f11;
    'h1096: romdata_int = 'h3000;
    'h1097: romdata_int = 'h650b;
    'h1098: romdata_int = 'h6e08;
    'h1099: romdata_int = 'h7800;
    'h109a: romdata_int = 'h9530;
    'h109b: romdata_int = 'hc000;
    'h109c: romdata_int = 'hcec5;
    'h109d: romdata_int = 'hdad7;
    'h109e: romdata_int = 'h10800;
    'h109f: romdata_int = 'h11230;
    'h10a0: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h10a1: romdata_int = 'h718;
    'h10a2: romdata_int = 'h1a16;
    'h10a3: romdata_int = 'h1c7d;
    'h10a4: romdata_int = 'h22d9;
    'h10a5: romdata_int = 'h234c;
    'h10a6: romdata_int = 'h3200;
    'h10a7: romdata_int = 'h3836;
    'h10a8: romdata_int = 'h7a00;
    'h10a9: romdata_int = 'h80cd;
    'h10aa: romdata_int = 'h8151;
    'h10ab: romdata_int = 'hbf12;
    'h10ac: romdata_int = 'hc200;
    'h10ad: romdata_int = 'hcd2f;
    'h10ae: romdata_int = 'hea87;
    'h10af: romdata_int = 'h10a00;
    'h10b0: romdata_int = 'h10a7b;
    'h10b1: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h10b2: romdata_int = 'h267;
    'h10b3: romdata_int = 'hc28;
    'h10b4: romdata_int = 'h1273;
    'h10b5: romdata_int = 'h14e4;
    'h10b6: romdata_int = 'h1a7a;
    'h10b7: romdata_int = 'h291c;
    'h10b8: romdata_int = 'h3400;
    'h10b9: romdata_int = 'h50b8;
    'h10ba: romdata_int = 'h64f4;
    'h10bb: romdata_int = 'h7c00;
    'h10bc: romdata_int = 'h94df;
    'h10bd: romdata_int = 'hae29;
    'h10be: romdata_int = 'hc400;
    'h10bf: romdata_int = 'he613;
    'h10c0: romdata_int = 'hef16;
    'h10c1: romdata_int = 'h10c00;
    'h10c2: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h10c3: romdata_int = 'hd38;
    'h10c4: romdata_int = 'h107b;
    'h10c5: romdata_int = 'h1282;
    'h10c6: romdata_int = 'h14f6;
    'h10c7: romdata_int = 'h1a28;
    'h10c8: romdata_int = 'h1e6f;
    'h10c9: romdata_int = 'h3600;
    'h10ca: romdata_int = 'h5932;
    'h10cb: romdata_int = 'h7e00;
    'h10cc: romdata_int = 'h847b;
    'h10cd: romdata_int = 'haaa7;
    'h10ce: romdata_int = 'hb4c2;
    'h10cf: romdata_int = 'hc600;
    'h10d0: romdata_int = 'h10e00;
    'h10d1: romdata_int = 'h118d0;
    'h10d2: romdata_int = 'h11c6f;
    'h10d3: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h10d4: romdata_int = 'h613;
    'h10d5: romdata_int = 'h6d0;
    'h10d6: romdata_int = 'hb2a;
    'h10d7: romdata_int = 'hc21;
    'h10d8: romdata_int = 'h22d4;
    'h10d9: romdata_int = 'h314c;
    'h10da: romdata_int = 'h3800;
    'h10db: romdata_int = 'h5243;
    'h10dc: romdata_int = 'h7553;
    'h10dd: romdata_int = 'h8000;
    'h10de: romdata_int = 'hba8d;
    'h10df: romdata_int = 'hc800;
    'h10e0: romdata_int = 'hcaf1;
    'h10e1: romdata_int = 'hf00b;
    'h10e2: romdata_int = 'h1046a;
    'h10e3: romdata_int = 'h11000;
    'h10e4: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h10e5: romdata_int = 'h4c4;
    'h10e6: romdata_int = 'h1907;
    'h10e7: romdata_int = 'h1a0e;
    'h10e8: romdata_int = 'h1c2a;
    'h10e9: romdata_int = 'h20db;
    'h10ea: romdata_int = 'h393e;
    'h10eb: romdata_int = 'h3a00;
    'h10ec: romdata_int = 'h6a22;
    'h10ed: romdata_int = 'h6ed2;
    'h10ee: romdata_int = 'h8200;
    'h10ef: romdata_int = 'hb21a;
    'h10f0: romdata_int = 'hc4b9;
    'h10f1: romdata_int = 'hca00;
    'h10f2: romdata_int = 'h11200;
    'h10f3: romdata_int = 'h1140d;
    'h10f4: romdata_int = 'h11d56;
    'h10f5: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h10f6: romdata_int = 'h28a;
    'h10f7: romdata_int = 'h4f2;
    'h10f8: romdata_int = 'h103e;
    'h10f9: romdata_int = 'h1c52;
    'h10fa: romdata_int = 'h2155;
    'h10fb: romdata_int = 'h3c00;
    'h10fc: romdata_int = 'h4752;
    'h10fd: romdata_int = 'h5f54;
    'h10fe: romdata_int = 'h6696;
    'h10ff: romdata_int = 'h8400;
    'h1100: romdata_int = 'hbcbf;
    'h1101: romdata_int = 'hcc00;
    'h1102: romdata_int = 'hd28e;
    'h1103: romdata_int = 'he011;
    'h1104: romdata_int = 'he415;
    'h1105: romdata_int = 'h11400;
    'h1106: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h1107: romdata_int = 'h9a;
    'h1108: romdata_int = 'h15c;
    'h1109: romdata_int = 'h10db;
    'h110a: romdata_int = 'h1a91;
    'h110b: romdata_int = 'h2f54;
    'h110c: romdata_int = 'h3e00;
    'h110d: romdata_int = 'h4562;
    'h110e: romdata_int = 'h4a9b;
    'h110f: romdata_int = 'h8600;
    'h1110: romdata_int = 'h8e6f;
    'h1111: romdata_int = 'h909c;
    'h1112: romdata_int = 'ha06b;
    'h1113: romdata_int = 'hce00;
    'h1114: romdata_int = 'hdb2d;
    'h1115: romdata_int = 'hdd56;
    'h1116: romdata_int = 'h11600;
    'h1117: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h1118: romdata_int = 'h255;
    'h1119: romdata_int = 'h10c3;
    'h111a: romdata_int = 'h1738;
    'h111b: romdata_int = 'h1d08;
    'h111c: romdata_int = 'h30bd;
    'h111d: romdata_int = 'h3efc;
    'h111e: romdata_int = 'h4000;
    'h111f: romdata_int = 'h568e;
    'h1120: romdata_int = 'h60d2;
    'h1121: romdata_int = 'h8800;
    'h1122: romdata_int = 'ha4a5;
    'h1123: romdata_int = 'hb646;
    'h1124: romdata_int = 'hd000;
    'h1125: romdata_int = 'h108f0;
    'h1126: romdata_int = 'h11800;
    'h1127: romdata_int = 'h11a4a;
    'h1128: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h1129: romdata_int = 'h43b;
    'h112a: romdata_int = 'h64e;
    'h112b: romdata_int = 'h80e;
    'h112c: romdata_int = 'h126b;
    'h112d: romdata_int = 'h191e;
    'h112e: romdata_int = 'h2030;
    'h112f: romdata_int = 'h4200;
    'h1130: romdata_int = 'h493d;
    'h1131: romdata_int = 'h8547;
    'h1132: romdata_int = 'h8a00;
    'h1133: romdata_int = 'hbe3a;
    'h1134: romdata_int = 'hceae;
    'h1135: romdata_int = 'hd200;
    'h1136: romdata_int = 'he453;
    'h1137: romdata_int = 'h11844;
    'h1138: romdata_int = 'h11a00;
    'h1139: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h113a: romdata_int = 'h6e7;
    'h113b: romdata_int = 'h875;
    'h113c: romdata_int = 'h1267;
    'h113d: romdata_int = 'h14dc;
    'h113e: romdata_int = 'h2474;
    'h113f: romdata_int = 'h40cb;
    'h1140: romdata_int = 'h4400;
    'h1141: romdata_int = 'h4acf;
    'h1142: romdata_int = 'h76f3;
    'h1143: romdata_int = 'h8c00;
    'h1144: romdata_int = 'h9233;
    'h1145: romdata_int = 'ha866;
    'h1146: romdata_int = 'hd400;
    'h1147: romdata_int = 'he639;
    'h1148: romdata_int = 'hfcbd;
    'h1149: romdata_int = 'h11c00;
    'h114a: romdata_int = 'h6f24; // Line descriptor for 4_5
    'h114b: romdata_int = 'h2d5;
    'h114c: romdata_int = 'h64a;
    'h114d: romdata_int = 'h938;
    'h114e: romdata_int = 'h14ef;
    'h114f: romdata_int = 'h1839;
    'h1150: romdata_int = 'h2e6b;
    'h1151: romdata_int = 'h4600;
    'h1152: romdata_int = 'h4c77;
    'h1153: romdata_int = 'h8e00;
    'h1154: romdata_int = 'h8e1f;
    'h1155: romdata_int = 'hb638;
    'h1156: romdata_int = 'hcce2;
    'h1157: romdata_int = 'hd600;
    'h1158: romdata_int = 'hd911;
    'h1159: romdata_int = 'h10f50;
    'h115a: romdata_int = 'h11e00;
    'h115b: romdata_int = 'h531e; // Line descriptor for 5_6
    'h115c: romdata_int = 'h0;
    'h115d: romdata_int = 'h738;
    'h115e: romdata_int = 'hd4c;
    'h115f: romdata_int = 'h1056;
    'h1160: romdata_int = 'h1280;
    'h1161: romdata_int = 'h1a8e;
    'h1162: romdata_int = 'h1c13;
    'h1163: romdata_int = 'h1c78;
    'h1164: romdata_int = 'h3c00;
    'h1165: romdata_int = 'h5058;
    'h1166: romdata_int = 'h6d18;
    'h1167: romdata_int = 'h7800;
    'h1168: romdata_int = 'h9118;
    'h1169: romdata_int = 'h9c15;
    'h116a: romdata_int = 'hb400;
    'h116b: romdata_int = 'hc26c;
    'h116c: romdata_int = 'heca1;
    'h116d: romdata_int = 'hf000;
    'h116e: romdata_int = 'h1106f;
    'h116f: romdata_int = 'h11897;
    'h1170: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1171: romdata_int = 'h200;
    'h1172: romdata_int = 'h2c9;
    'h1173: romdata_int = 'h467;
    'h1174: romdata_int = 'h4bd;
    'h1175: romdata_int = 'hf07;
    'h1176: romdata_int = 'h1adf;
    'h1177: romdata_int = 'h1efe;
    'h1178: romdata_int = 'h271c;
    'h1179: romdata_int = 'h3e00;
    'h117a: romdata_int = 'h3e58;
    'h117b: romdata_int = 'h5d11;
    'h117c: romdata_int = 'h7a00;
    'h117d: romdata_int = 'h86ab;
    'h117e: romdata_int = 'h8ad3;
    'h117f: romdata_int = 'hb600;
    'h1180: romdata_int = 'hc8bf;
    'h1181: romdata_int = 'hcacc;
    'h1182: romdata_int = 'hf200;
    'h1183: romdata_int = 'h1062b;
    'h1184: romdata_int = 'h12847;
    'h1185: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1186: romdata_int = 'h61;
    'h1187: romdata_int = 'h400;
    'h1188: romdata_int = 'ha87;
    'h1189: romdata_int = 'h12db;
    'h118a: romdata_int = 'h18f5;
    'h118b: romdata_int = 'h193e;
    'h118c: romdata_int = 'h36a9;
    'h118d: romdata_int = 'h3876;
    'h118e: romdata_int = 'h4000;
    'h118f: romdata_int = 'h54ba;
    'h1190: romdata_int = 'h70a8;
    'h1191: romdata_int = 'h7c00;
    'h1192: romdata_int = 'h829b;
    'h1193: romdata_int = 'h8cde;
    'h1194: romdata_int = 'hb678;
    'h1195: romdata_int = 'hb800;
    'h1196: romdata_int = 'he80c;
    'h1197: romdata_int = 'hf400;
    'h1198: romdata_int = 'h104cc;
    'h1199: romdata_int = 'h10961;
    'h119a: romdata_int = 'h531e; // Line descriptor for 5_6
    'h119b: romdata_int = 'he0;
    'h119c: romdata_int = 'h600;
    'h119d: romdata_int = 'h948;
    'h119e: romdata_int = 'ha7b;
    'h119f: romdata_int = 'h1060;
    'h11a0: romdata_int = 'h1761;
    'h11a1: romdata_int = 'h1962;
    'h11a2: romdata_int = 'h22f3;
    'h11a3: romdata_int = 'h4200;
    'h11a4: romdata_int = 'h44fa;
    'h11a5: romdata_int = 'h74f0;
    'h11a6: romdata_int = 'h7e00;
    'h11a7: romdata_int = 'h80d9;
    'h11a8: romdata_int = 'h9e0c;
    'h11a9: romdata_int = 'hb469;
    'h11aa: romdata_int = 'hba00;
    'h11ab: romdata_int = 'hde19;
    'h11ac: romdata_int = 'hf600;
    'h11ad: romdata_int = 'h11360;
    'h11ae: romdata_int = 'h1289c;
    'h11af: romdata_int = 'h531e; // Line descriptor for 5_6
    'h11b0: romdata_int = 'h800;
    'h11b1: romdata_int = 'h905;
    'h11b2: romdata_int = 'haee;
    'h11b3: romdata_int = 'h1022;
    'h11b4: romdata_int = 'h1245;
    'h11b5: romdata_int = 'h1267;
    'h11b6: romdata_int = 'h160d;
    'h11b7: romdata_int = 'h1ed2;
    'h11b8: romdata_int = 'h4400;
    'h11b9: romdata_int = 'h4e84;
    'h11ba: romdata_int = 'h6e0d;
    'h11bb: romdata_int = 'h8000;
    'h11bc: romdata_int = 'h9a5f;
    'h11bd: romdata_int = 'haeca;
    'h11be: romdata_int = 'hbc00;
    'h11bf: romdata_int = 'hdb2e;
    'h11c0: romdata_int = 'he257;
    'h11c1: romdata_int = 'hf800;
    'h11c2: romdata_int = 'h1128e;
    'h11c3: romdata_int = 'h124d6;
    'h11c4: romdata_int = 'h531e; // Line descriptor for 5_6
    'h11c5: romdata_int = 'h4a6;
    'h11c6: romdata_int = 'h553;
    'h11c7: romdata_int = 'h8a1;
    'h11c8: romdata_int = 'ha00;
    'h11c9: romdata_int = 'he9e;
    'h11ca: romdata_int = 'h1049;
    'h11cb: romdata_int = 'h1818;
    'h11cc: romdata_int = 'h1a7d;
    'h11cd: romdata_int = 'h4600;
    'h11ce: romdata_int = 'h606e;
    'h11cf: romdata_int = 'h6f13;
    'h11d0: romdata_int = 'h7f61;
    'h11d1: romdata_int = 'h8200;
    'h11d2: romdata_int = 'hb260;
    'h11d3: romdata_int = 'hb687;
    'h11d4: romdata_int = 'hbe00;
    'h11d5: romdata_int = 'he645;
    'h11d6: romdata_int = 'hfa00;
    'h11d7: romdata_int = 'h1092a;
    'h11d8: romdata_int = 'h1267d;
    'h11d9: romdata_int = 'h531e; // Line descriptor for 5_6
    'h11da: romdata_int = 'h6b;
    'h11db: romdata_int = 'h74d;
    'h11dc: romdata_int = 'hc00;
    'h11dd: romdata_int = 'hd15;
    'h11de: romdata_int = 'he8b;
    'h11df: romdata_int = 'h127e;
    'h11e0: romdata_int = 'h1679;
    'h11e1: romdata_int = 'h22e2;
    'h11e2: romdata_int = 'h4800;
    'h11e3: romdata_int = 'h4b35;
    'h11e4: romdata_int = 'h5a96;
    'h11e5: romdata_int = 'h8400;
    'h11e6: romdata_int = 'h9331;
    'h11e7: romdata_int = 'hac97;
    'h11e8: romdata_int = 'hc000;
    'h11e9: romdata_int = 'hd70b;
    'h11ea: romdata_int = 'hdef4;
    'h11eb: romdata_int = 'hfc00;
    'h11ec: romdata_int = 'h10342;
    'h11ed: romdata_int = 'h11e46;
    'h11ee: romdata_int = 'h531e; // Line descriptor for 5_6
    'h11ef: romdata_int = 'h2d5;
    'h11f0: romdata_int = 'h4f2;
    'h11f1: romdata_int = 'h68f;
    'h11f2: romdata_int = 'he34;
    'h11f3: romdata_int = 'he00;
    'h11f4: romdata_int = 'he39;
    'h11f5: romdata_int = 'h2d3d;
    'h11f6: romdata_int = 'h3623;
    'h11f7: romdata_int = 'h4a00;
    'h11f8: romdata_int = 'h5ecd;
    'h11f9: romdata_int = 'h6825;
    'h11fa: romdata_int = 'h7c02;
    'h11fb: romdata_int = 'h8600;
    'h11fc: romdata_int = 'ha6c0;
    'h11fd: romdata_int = 'hb839;
    'h11fe: romdata_int = 'hc200;
    'h11ff: romdata_int = 'he89c;
    'h1200: romdata_int = 'hf105;
    'h1201: romdata_int = 'hf67a;
    'h1202: romdata_int = 'hfe00;
    'h1203: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1204: romdata_int = 'h32b;
    'h1205: romdata_int = 'h6ab;
    'h1206: romdata_int = 'h74f;
    'h1207: romdata_int = 'h1000;
    'h1208: romdata_int = 'h18fc;
    'h1209: romdata_int = 'h1b25;
    'h120a: romdata_int = 'h2d56;
    'h120b: romdata_int = 'h3908;
    'h120c: romdata_int = 'h4c00;
    'h120d: romdata_int = 'h4e0b;
    'h120e: romdata_int = 'h70d3;
    'h120f: romdata_int = 'h7cf1;
    'h1210: romdata_int = 'h8800;
    'h1211: romdata_int = 'h8f55;
    'h1212: romdata_int = 'hbd07;
    'h1213: romdata_int = 'hc400;
    'h1214: romdata_int = 'hc906;
    'h1215: romdata_int = 'h10000;
    'h1216: romdata_int = 'h104ec;
    'h1217: romdata_int = 'h11ae3;
    'h1218: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1219: romdata_int = 'h52c;
    'h121a: romdata_int = 'h84f;
    'h121b: romdata_int = 'hc17;
    'h121c: romdata_int = 'hcad;
    'h121d: romdata_int = 'h1038;
    'h121e: romdata_int = 'h1094;
    'h121f: romdata_int = 'h1200;
    'h1220: romdata_int = 'h1af7;
    'h1221: romdata_int = 'h4e00;
    'h1222: romdata_int = 'h6abb;
    'h1223: romdata_int = 'h7442;
    'h1224: romdata_int = 'h8a00;
    'h1225: romdata_int = 'h9b1a;
    'h1226: romdata_int = 'ha52e;
    'h1227: romdata_int = 'hc53c;
    'h1228: romdata_int = 'hc600;
    'h1229: romdata_int = 'hd264;
    'h122a: romdata_int = 'hf238;
    'h122b: romdata_int = 'h10200;
    'h122c: romdata_int = 'h10a78;
    'h122d: romdata_int = 'h531e; // Line descriptor for 5_6
    'h122e: romdata_int = 'h55;
    'h122f: romdata_int = 'h670;
    'h1230: romdata_int = 'h866;
    'h1231: romdata_int = 'h1230;
    'h1232: romdata_int = 'h1400;
    'h1233: romdata_int = 'h1cd9;
    'h1234: romdata_int = 'h24c6;
    'h1235: romdata_int = 'h30b9;
    'h1236: romdata_int = 'h4539;
    'h1237: romdata_int = 'h5000;
    'h1238: romdata_int = 'h6233;
    'h1239: romdata_int = 'h8c00;
    'h123a: romdata_int = 'h9838;
    'h123b: romdata_int = 'ha687;
    'h123c: romdata_int = 'hc800;
    'h123d: romdata_int = 'hce13;
    'h123e: romdata_int = 'heb4b;
    'h123f: romdata_int = 'h1006e;
    'h1240: romdata_int = 'h10400;
    'h1241: romdata_int = 'h10aed;
    'h1242: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1243: romdata_int = 'h264;
    'h1244: romdata_int = 'hb06;
    'h1245: romdata_int = 'hc42;
    'h1246: romdata_int = 'hd58;
    'h1247: romdata_int = 'h1600;
    'h1248: romdata_int = 'h171d;
    'h1249: romdata_int = 'h1854;
    'h124a: romdata_int = 'h1aee;
    'h124b: romdata_int = 'h5200;
    'h124c: romdata_int = 'h5a74;
    'h124d: romdata_int = 'h763b;
    'h124e: romdata_int = 'h7f26;
    'h124f: romdata_int = 'h8e00;
    'h1250: romdata_int = 'hb244;
    'h1251: romdata_int = 'hb564;
    'h1252: romdata_int = 'hca00;
    'h1253: romdata_int = 'he614;
    'h1254: romdata_int = 'h10600;
    'h1255: romdata_int = 'h120e5;
    'h1256: romdata_int = 'h12248;
    'h1257: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1258: romdata_int = 'h91;
    'h1259: romdata_int = 'h488;
    'h125a: romdata_int = 'hf66;
    'h125b: romdata_int = 'h1232;
    'h125c: romdata_int = 'h153b;
    'h125d: romdata_int = 'h1681;
    'h125e: romdata_int = 'h1800;
    'h125f: romdata_int = 'h3a7d;
    'h1260: romdata_int = 'h4a38;
    'h1261: romdata_int = 'h5400;
    'h1262: romdata_int = 'h5c8b;
    'h1263: romdata_int = 'h9000;
    'h1264: romdata_int = 'ha2df;
    'h1265: romdata_int = 'had28;
    'h1266: romdata_int = 'hc4de;
    'h1267: romdata_int = 'hcc00;
    'h1268: romdata_int = 'hcd30;
    'h1269: romdata_int = 'h10800;
    'h126a: romdata_int = 'h10f0c;
    'h126b: romdata_int = 'h12487;
    'h126c: romdata_int = 'h531e; // Line descriptor for 5_6
    'h126d: romdata_int = 'h11e;
    'h126e: romdata_int = 'h336;
    'h126f: romdata_int = 'h916;
    'h1270: romdata_int = 'hee5;
    'h1271: romdata_int = 'h131e;
    'h1272: romdata_int = 'h1836;
    'h1273: romdata_int = 'h1a00;
    'h1274: romdata_int = 'h1b13;
    'h1275: romdata_int = 'h54bd;
    'h1276: romdata_int = 'h5600;
    'h1277: romdata_int = 'h573d;
    'h1278: romdata_int = 'h9200;
    'h1279: romdata_int = 'hae1c;
    'h127a: romdata_int = 'hb0c4;
    'h127b: romdata_int = 'hcca1;
    'h127c: romdata_int = 'hce00;
    'h127d: romdata_int = 'hee2d;
    'h127e: romdata_int = 'h10a00;
    'h127f: romdata_int = 'h11c71;
    'h1280: romdata_int = 'h12081;
    'h1281: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1282: romdata_int = 'h60e;
    'h1283: romdata_int = 'ha45;
    'h1284: romdata_int = 'hc2b;
    'h1285: romdata_int = 'hf45;
    'h1286: romdata_int = 'h12b5;
    'h1287: romdata_int = 'h1711;
    'h1288: romdata_int = 'h1802;
    'h1289: romdata_int = 'h1c00;
    'h128a: romdata_int = 'h405c;
    'h128b: romdata_int = 'h5800;
    'h128c: romdata_int = 'h76ac;
    'h128d: romdata_int = 'h7a8c;
    'h128e: romdata_int = 'h8f40;
    'h128f: romdata_int = 'h9400;
    'h1290: romdata_int = 'hd000;
    'h1291: romdata_int = 'he305;
    'h1292: romdata_int = 'heb21;
    'h1293: romdata_int = 'hfa8d;
    'h1294: romdata_int = 'hfe83;
    'h1295: romdata_int = 'h10c00;
    'h1296: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1297: romdata_int = 'hd5;
    'h1298: romdata_int = 'ha72;
    'h1299: romdata_int = 'hadb;
    'h129a: romdata_int = 'h154c;
    'h129b: romdata_int = 'h1708;
    'h129c: romdata_int = 'h1c42;
    'h129d: romdata_int = 'h1e00;
    'h129e: romdata_int = 'h3212;
    'h129f: romdata_int = 'h3f41;
    'h12a0: romdata_int = 'h5a00;
    'h12a1: romdata_int = 'h66de;
    'h12a2: romdata_int = 'h910b;
    'h12a3: romdata_int = 'h9600;
    'h12a4: romdata_int = 'ha089;
    'h12a5: romdata_int = 'hd200;
    'h12a6: romdata_int = 'hd406;
    'h12a7: romdata_int = 'hd932;
    'h12a8: romdata_int = 'hfd55;
    'h12a9: romdata_int = 'h10e00;
    'h12aa: romdata_int = 'h11060;
    'h12ab: romdata_int = 'h531e; // Line descriptor for 5_6
    'h12ac: romdata_int = 'h8a;
    'h12ad: romdata_int = 'h23b;
    'h12ae: romdata_int = 'h522;
    'h12af: romdata_int = 'ha3e;
    'h12b0: romdata_int = 'h10d8;
    'h12b1: romdata_int = 'h1cb5;
    'h12b2: romdata_int = 'h2000;
    'h12b3: romdata_int = 'h3a6b;
    'h12b4: romdata_int = 'h495c;
    'h12b5: romdata_int = 'h561e;
    'h12b6: romdata_int = 'h5c00;
    'h12b7: romdata_int = 'h7a70;
    'h12b8: romdata_int = 'h9800;
    'h12b9: romdata_int = 'ha533;
    'h12ba: romdata_int = 'hd400;
    'h12bb: romdata_int = 'hd832;
    'h12bc: romdata_int = 'he415;
    'h12bd: romdata_int = 'h102d3;
    'h12be: romdata_int = 'h11000;
    'h12bf: romdata_int = 'h114d8;
    'h12c0: romdata_int = 'h531e; // Line descriptor for 5_6
    'h12c1: romdata_int = 'h262;
    'h12c2: romdata_int = 'h354;
    'h12c3: romdata_int = 'h45c;
    'h12c4: romdata_int = 'h84d;
    'h12c5: romdata_int = 'hc82;
    'h12c6: romdata_int = 'h12a8;
    'h12c7: romdata_int = 'h2200;
    'h12c8: romdata_int = 'h347f;
    'h12c9: romdata_int = 'h4d4e;
    'h12ca: romdata_int = 'h50a9;
    'h12cb: romdata_int = 'h5e00;
    'h12cc: romdata_int = 'h8ab7;
    'h12cd: romdata_int = 'h94eb;
    'h12ce: romdata_int = 'h9a00;
    'h12cf: romdata_int = 'hbe14;
    'h12d0: romdata_int = 'hc6f8;
    'h12d1: romdata_int = 'hd600;
    'h12d2: romdata_int = 'h11200;
    'h12d3: romdata_int = 'h11725;
    'h12d4: romdata_int = 'h12b0b;
    'h12d5: romdata_int = 'h531e; // Line descriptor for 5_6
    'h12d6: romdata_int = 'h625;
    'h12d7: romdata_int = 'ha0b;
    'h12d8: romdata_int = 'he81;
    'h12d9: romdata_int = 'h143d;
    'h12da: romdata_int = 'h174c;
    'h12db: romdata_int = 'h1c19;
    'h12dc: romdata_int = 'h20d8;
    'h12dd: romdata_int = 'h2400;
    'h12de: romdata_int = 'h4c86;
    'h12df: romdata_int = 'h521c;
    'h12e0: romdata_int = 'h6000;
    'h12e1: romdata_int = 'h8706;
    'h12e2: romdata_int = 'h9c00;
    'h12e3: romdata_int = 'ha0e9;
    'h12e4: romdata_int = 'hd24b;
    'h12e5: romdata_int = 'hd800;
    'h12e6: romdata_int = 'heeea;
    'h12e7: romdata_int = 'hf74a;
    'h12e8: romdata_int = 'h10d31;
    'h12e9: romdata_int = 'h11400;
    'h12ea: romdata_int = 'h531e; // Line descriptor for 5_6
    'h12eb: romdata_int = 'ha5;
    'h12ec: romdata_int = 'h252;
    'h12ed: romdata_int = 'h290;
    'h12ee: romdata_int = 'h549;
    'h12ef: romdata_int = 'hf4d;
    'h12f0: romdata_int = 'h14d4;
    'h12f1: romdata_int = 'h2600;
    'h12f2: romdata_int = 'h2f37;
    'h12f3: romdata_int = 'h6200;
    'h12f4: romdata_int = 'h6687;
    'h12f5: romdata_int = 'h72aa;
    'h12f6: romdata_int = 'h7876;
    'h12f7: romdata_int = 'h842f;
    'h12f8: romdata_int = 'h9e00;
    'h12f9: romdata_int = 'hbc40;
    'h12fa: romdata_int = 'hd450;
    'h12fb: romdata_int = 'hda00;
    'h12fc: romdata_int = 'hf44e;
    'h12fd: romdata_int = 'h11600;
    'h12fe: romdata_int = 'h11842;
    'h12ff: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1300: romdata_int = 'hac3;
    'h1301: romdata_int = 'ha5c;
    'h1302: romdata_int = 'hb58;
    'h1303: romdata_int = 'h10b4;
    'h1304: romdata_int = 'h1c06;
    'h1305: romdata_int = 'h2800;
    'h1306: romdata_int = 'h2a27;
    'h1307: romdata_int = 'h351e;
    'h1308: romdata_int = 'h3c50;
    'h1309: romdata_int = 'h463d;
    'h130a: romdata_int = 'h6400;
    'h130b: romdata_int = 'h82b0;
    'h130c: romdata_int = 'h92bb;
    'h130d: romdata_int = 'ha000;
    'h130e: romdata_int = 'hc669;
    'h130f: romdata_int = 'hd135;
    'h1310: romdata_int = 'hdc00;
    'h1311: romdata_int = 'hf54f;
    'h1312: romdata_int = 'hf8e6;
    'h1313: romdata_int = 'h11800;
    'h1314: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1315: romdata_int = 'h8f3;
    'h1316: romdata_int = 'hc35;
    'h1317: romdata_int = 'hc67;
    'h1318: romdata_int = 'h1003;
    'h1319: romdata_int = 'h126e;
    'h131a: romdata_int = 'h1ce1;
    'h131b: romdata_int = 'h2a00;
    'h131c: romdata_int = 'h2e48;
    'h131d: romdata_int = 'h4243;
    'h131e: romdata_int = 'h42b1;
    'h131f: romdata_int = 'h6600;
    'h1320: romdata_int = 'h8028;
    'h1321: romdata_int = 'h8ca4;
    'h1322: romdata_int = 'ha200;
    'h1323: romdata_int = 'hcf3f;
    'h1324: romdata_int = 'hde00;
    'h1325: romdata_int = 'he0d1;
    'h1326: romdata_int = 'hf27e;
    'h1327: romdata_int = 'hfd04;
    'h1328: romdata_int = 'h11a00;
    'h1329: romdata_int = 'h531e; // Line descriptor for 5_6
    'h132a: romdata_int = 'h67;
    'h132b: romdata_int = 'h72d;
    'h132c: romdata_int = 'h1349;
    'h132d: romdata_int = 'h1559;
    'h132e: romdata_int = 'h1a45;
    'h132f: romdata_int = 'h1a52;
    'h1330: romdata_int = 'h1d28;
    'h1331: romdata_int = 'h2c00;
    'h1332: romdata_int = 'h4051;
    'h1333: romdata_int = 'h5f53;
    'h1334: romdata_int = 'h6800;
    'h1335: romdata_int = 'ha235;
    'h1336: romdata_int = 'ha400;
    'h1337: romdata_int = 'haab9;
    'h1338: romdata_int = 'hcb65;
    'h1339: romdata_int = 'hdb0c;
    'h133a: romdata_int = 'he000;
    'h133b: romdata_int = 'h10d2f;
    'h133c: romdata_int = 'h11b32;
    'h133d: romdata_int = 'h11c00;
    'h133e: romdata_int = 'h531e; // Line descriptor for 5_6
    'h133f: romdata_int = 'h10c8;
    'h1340: romdata_int = 'h14f3;
    'h1341: romdata_int = 'h1aa6;
    'h1342: romdata_int = 'h1b32;
    'h1343: romdata_int = 'h1c24;
    'h1344: romdata_int = 'h263b;
    'h1345: romdata_int = 'h2b45;
    'h1346: romdata_int = 'h2e00;
    'h1347: romdata_int = 'h5273;
    'h1348: romdata_int = 'h6a00;
    'h1349: romdata_int = 'h6d1a;
    'h134a: romdata_int = 'h9eb5;
    'h134b: romdata_int = 'ha600;
    'h134c: romdata_int = 'ha87c;
    'h134d: romdata_int = 'he07f;
    'h134e: romdata_int = 'he200;
    'h134f: romdata_int = 'he44c;
    'h1350: romdata_int = 'h10ece;
    'h1351: romdata_int = 'h11e00;
    'h1352: romdata_int = 'h11f2c;
    'h1353: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1354: romdata_int = 'h2b6;
    'h1355: romdata_int = 'h527;
    'h1356: romdata_int = 'h682;
    'h1357: romdata_int = 'h81a;
    'h1358: romdata_int = 'he99;
    'h1359: romdata_int = 'h28cd;
    'h135a: romdata_int = 'h2905;
    'h135b: romdata_int = 'h3000;
    'h135c: romdata_int = 'h4945;
    'h135d: romdata_int = 'h6c00;
    'h135e: romdata_int = 'h72cd;
    'h135f: romdata_int = 'h7830;
    'h1360: romdata_int = 'h8956;
    'h1361: romdata_int = 'ha800;
    'h1362: romdata_int = 'hc02d;
    'h1363: romdata_int = 'hc11c;
    'h1364: romdata_int = 'he400;
    'h1365: romdata_int = 'hf83f;
    'h1366: romdata_int = 'h11c39;
    'h1367: romdata_int = 'h12000;
    'h1368: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1369: romdata_int = 'h69f;
    'h136a: romdata_int = 'h752;
    'h136b: romdata_int = 'h1498;
    'h136c: romdata_int = 'h164f;
    'h136d: romdata_int = 'h1903;
    'h136e: romdata_int = 'h192f;
    'h136f: romdata_int = 'h1b50;
    'h1370: romdata_int = 'h3200;
    'h1371: romdata_int = 'h3cea;
    'h1372: romdata_int = 'h6a66;
    'h1373: romdata_int = 'h6e00;
    'h1374: romdata_int = 'h8893;
    'h1375: romdata_int = 'h9671;
    'h1376: romdata_int = 'haa00;
    'h1377: romdata_int = 'hdc45;
    'h1378: romdata_int = 'he600;
    'h1379: romdata_int = 'hec44;
    'h137a: romdata_int = 'h116fe;
    'h137b: romdata_int = 'h12200;
    'h137c: romdata_int = 'h12281;
    'h137d: romdata_int = 'h531e; // Line descriptor for 5_6
    'h137e: romdata_int = 'hd;
    'h137f: romdata_int = 'hc73;
    'h1380: romdata_int = 'h143a;
    'h1381: romdata_int = 'h14ba;
    'h1382: romdata_int = 'h1451;
    'h1383: romdata_int = 'h14d9;
    'h1384: romdata_int = 'h3233;
    'h1385: romdata_int = 'h3400;
    'h1386: romdata_int = 'h649e;
    'h1387: romdata_int = 'h6821;
    'h1388: romdata_int = 'h7000;
    'h1389: romdata_int = 'h9880;
    'h138a: romdata_int = 'h9cce;
    'h138b: romdata_int = 'hac00;
    'h138c: romdata_int = 'hbe06;
    'h138d: romdata_int = 'hc363;
    'h138e: romdata_int = 'he800;
    'h138f: romdata_int = 'h1155f;
    'h1390: romdata_int = 'h12400;
    'h1391: romdata_int = 'h1273d;
    'h1392: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1393: romdata_int = 'h8ee;
    'h1394: romdata_int = 'he6b;
    'h1395: romdata_int = 'h1160;
    'h1396: romdata_int = 'h1734;
    'h1397: romdata_int = 'h18d5;
    'h1398: romdata_int = 'h18e4;
    'h1399: romdata_int = 'h1c96;
    'h139a: romdata_int = 'h3600;
    'h139b: romdata_int = 'h5888;
    'h139c: romdata_int = 'h6459;
    'h139d: romdata_int = 'h7200;
    'h139e: romdata_int = 'h972c;
    'h139f: romdata_int = 'ha933;
    'h13a0: romdata_int = 'hae00;
    'h13a1: romdata_int = 'hd0d0;
    'h13a2: romdata_int = 'hd633;
    'h13a3: romdata_int = 'hea00;
    'h13a4: romdata_int = 'h10704;
    'h13a5: romdata_int = 'h12600;
    'h13a6: romdata_int = 'h12af4;
    'h13a7: romdata_int = 'h531e; // Line descriptor for 5_6
    'h13a8: romdata_int = 'h2f2;
    'h13a9: romdata_int = 'h832;
    'h13aa: romdata_int = 'h1062;
    'h13ab: romdata_int = 'h151c;
    'h13ac: romdata_int = 'h16c6;
    'h13ad: romdata_int = 'h1d43;
    'h13ae: romdata_int = 'h2438;
    'h13af: romdata_int = 'h3800;
    'h13b0: romdata_int = 'h464d;
    'h13b1: romdata_int = 'h60bc;
    'h13b2: romdata_int = 'h7400;
    'h13b3: romdata_int = 'h9527;
    'h13b4: romdata_int = 'haae9;
    'h13b5: romdata_int = 'hb000;
    'h13b6: romdata_int = 'hb80a;
    'h13b7: romdata_int = 'hdd2a;
    'h13b8: romdata_int = 'hec00;
    'h13b9: romdata_int = 'hfefe;
    'h13ba: romdata_int = 'h100b6;
    'h13bb: romdata_int = 'h12800;
    'h13bc: romdata_int = 'h731e; // Line descriptor for 5_6
    'h13bd: romdata_int = 'h128;
    'h13be: romdata_int = 'h448;
    'h13bf: romdata_int = 'h80a;
    'h13c0: romdata_int = 'hcc5;
    'h13c1: romdata_int = 'h16f2;
    'h13c2: romdata_int = 'h2132;
    'h13c3: romdata_int = 'h3040;
    'h13c4: romdata_int = 'h3a00;
    'h13c5: romdata_int = 'h5833;
    'h13c6: romdata_int = 'h6272;
    'h13c7: romdata_int = 'h7600;
    'h13c8: romdata_int = 'h8544;
    'h13c9: romdata_int = 'hb10c;
    'h13ca: romdata_int = 'hb200;
    'h13cb: romdata_int = 'hba49;
    'h13cc: romdata_int = 'hbb35;
    'h13cd: romdata_int = 'hee00;
    'h13ce: romdata_int = 'hf03a;
    'h13cf: romdata_int = 'hfabc;
    'h13d0: romdata_int = 'h12a00;
    'h13d1: romdata_int = 'h5814; // Line descriptor for 8_9
    'h13d2: romdata_int = 'h0;
    'h13d3: romdata_int = 'h322;
    'h13d4: romdata_int = 'h1ec4;
    'h13d5: romdata_int = 'h22e7;
    'h13d6: romdata_int = 'h2800;
    'h13d7: romdata_int = 'h3338;
    'h13d8: romdata_int = 'h4479;
    'h13d9: romdata_int = 'h5000;
    'h13da: romdata_int = 'h6425;
    'h13db: romdata_int = 'h72ee;
    'h13dc: romdata_int = 'h7800;
    'h13dd: romdata_int = 'h9a1e;
    'h13de: romdata_int = 'h9e3f;
    'h13df: romdata_int = 'ha000;
    'h13e0: romdata_int = 'ha616;
    'h13e1: romdata_int = 'hb750;
    'h13e2: romdata_int = 'hc800;
    'h13e3: romdata_int = 'hdace;
    'h13e4: romdata_int = 'hdad6;
    'h13e5: romdata_int = 'hf000;
    'h13e6: romdata_int = 'hf35c;
    'h13e7: romdata_int = 'h110d8;
    'h13e8: romdata_int = 'h11800;
    'h13e9: romdata_int = 'h13050;
    'h13ea: romdata_int = 'h13222;
    'h13eb: romdata_int = 'h5814; // Line descriptor for 8_9
    'h13ec: romdata_int = 'h200;
    'h13ed: romdata_int = 'h75c;
    'h13ee: romdata_int = 'h10bc;
    'h13ef: romdata_int = 'h2277;
    'h13f0: romdata_int = 'h2a00;
    'h13f1: romdata_int = 'h3d48;
    'h13f2: romdata_int = 'h4631;
    'h13f3: romdata_int = 'h5200;
    'h13f4: romdata_int = 'h5650;
    'h13f5: romdata_int = 'h7733;
    'h13f6: romdata_int = 'h7a00;
    'h13f7: romdata_int = 'h7e35;
    'h13f8: romdata_int = 'h8523;
    'h13f9: romdata_int = 'ha200;
    'h13fa: romdata_int = 'hac4a;
    'h13fb: romdata_int = 'hb8e2;
    'h13fc: romdata_int = 'hca00;
    'h13fd: romdata_int = 'hd870;
    'h13fe: romdata_int = 'he74a;
    'h13ff: romdata_int = 'hf200;
    'h1400: romdata_int = 'h11132;
    'h1401: romdata_int = 'h112c6;
    'h1402: romdata_int = 'h11a00;
    'h1403: romdata_int = 'h1345a;
    'h1404: romdata_int = 'h13854;
    'h1405: romdata_int = 'h5814; // Line descriptor for 8_9
    'h1406: romdata_int = 'ha1;
    'h1407: romdata_int = 'h400;
    'h1408: romdata_int = 'hf3d;
    'h1409: romdata_int = 'h224a;
    'h140a: romdata_int = 'h2c00;
    'h140b: romdata_int = 'h3b05;
    'h140c: romdata_int = 'h4cbe;
    'h140d: romdata_int = 'h5400;
    'h140e: romdata_int = 'h5719;
    'h140f: romdata_int = 'h6eeb;
    'h1410: romdata_int = 'h7c00;
    'h1411: romdata_int = 'h915d;
    'h1412: romdata_int = 'h98f2;
    'h1413: romdata_int = 'ha400;
    'h1414: romdata_int = 'hb6b5;
    'h1415: romdata_int = 'hc458;
    'h1416: romdata_int = 'hca67;
    'h1417: romdata_int = 'hcc00;
    'h1418: romdata_int = 'hd276;
    'h1419: romdata_int = 'hf400;
    'h141a: romdata_int = 'hf561;
    'h141b: romdata_int = 'h1007b;
    'h141c: romdata_int = 'h11c00;
    'h141d: romdata_int = 'h12904;
    'h141e: romdata_int = 'h12aec;
    'h141f: romdata_int = 'h5814; // Line descriptor for 8_9
    'h1420: romdata_int = 'h600;
    'h1421: romdata_int = 'hab8;
    'h1422: romdata_int = 'h1a43;
    'h1423: romdata_int = 'h1b28;
    'h1424: romdata_int = 'h2e00;
    'h1425: romdata_int = 'h3475;
    'h1426: romdata_int = 'h48d0;
    'h1427: romdata_int = 'h5600;
    'h1428: romdata_int = 'h5b21;
    'h1429: romdata_int = 'h6a70;
    'h142a: romdata_int = 'h7e00;
    'h142b: romdata_int = 'h7ead;
    'h142c: romdata_int = 'h9ef5;
    'h142d: romdata_int = 'ha41d;
    'h142e: romdata_int = 'ha600;
    'h142f: romdata_int = 'hb4c8;
    'h1430: romdata_int = 'hce00;
    'h1431: romdata_int = 'he446;
    'h1432: romdata_int = 'he703;
    'h1433: romdata_int = 'hf600;
    'h1434: romdata_int = 'h10738;
    'h1435: romdata_int = 'h10cad;
    'h1436: romdata_int = 'h11e00;
    'h1437: romdata_int = 'h122ca;
    'h1438: romdata_int = 'h1387b;
    'h1439: romdata_int = 'h5814; // Line descriptor for 8_9
    'h143a: romdata_int = 'h800;
    'h143b: romdata_int = 'h939;
    'h143c: romdata_int = 'h120d;
    'h143d: romdata_int = 'h2052;
    'h143e: romdata_int = 'h2a4b;
    'h143f: romdata_int = 'h2c5f;
    'h1440: romdata_int = 'h3000;
    'h1441: romdata_int = 'h5800;
    'h1442: romdata_int = 'h581a;
    'h1443: romdata_int = 'h6693;
    'h1444: romdata_int = 'h8000;
    'h1445: romdata_int = 'h8eb3;
    'h1446: romdata_int = 'h94f8;
    'h1447: romdata_int = 'ha2a1;
    'h1448: romdata_int = 'ha800;
    'h1449: romdata_int = 'hba3a;
    'h144a: romdata_int = 'hd000;
    'h144b: romdata_int = 'hed35;
    'h144c: romdata_int = 'hef52;
    'h144d: romdata_int = 'hf6b4;
    'h144e: romdata_int = 'hf800;
    'h144f: romdata_int = 'h10884;
    'h1450: romdata_int = 'h12000;
    'h1451: romdata_int = 'h12a97;
    'h1452: romdata_int = 'h13cd6;
    'h1453: romdata_int = 'h5814; // Line descriptor for 8_9
    'h1454: romdata_int = 'ha00;
    'h1455: romdata_int = 'ha79;
    'h1456: romdata_int = 'h18f3;
    'h1457: romdata_int = 'h192c;
    'h1458: romdata_int = 'h3200;
    'h1459: romdata_int = 'h3711;
    'h145a: romdata_int = 'h3eee;
    'h145b: romdata_int = 'h592c;
    'h145c: romdata_int = 'h5a00;
    'h145d: romdata_int = 'h7072;
    'h145e: romdata_int = 'h7a07;
    'h145f: romdata_int = 'h8200;
    'h1460: romdata_int = 'h98f6;
    'h1461: romdata_int = 'haa00;
    'h1462: romdata_int = 'hb267;
    'h1463: romdata_int = 'hbc62;
    'h1464: romdata_int = 'hd200;
    'h1465: romdata_int = 'hdd23;
    'h1466: romdata_int = 'he410;
    'h1467: romdata_int = 'hfa00;
    'h1468: romdata_int = 'hfe7d;
    'h1469: romdata_int = 'h11238;
    'h146a: romdata_int = 'h120c2;
    'h146b: romdata_int = 'h12200;
    'h146c: romdata_int = 'h12d10;
    'h146d: romdata_int = 'h5814; // Line descriptor for 8_9
    'h146e: romdata_int = 'hc00;
    'h146f: romdata_int = 'h1291;
    'h1470: romdata_int = 'h18a4;
    'h1471: romdata_int = 'h26bd;
    'h1472: romdata_int = 'h2934;
    'h1473: romdata_int = 'h3400;
    'h1474: romdata_int = 'h412a;
    'h1475: romdata_int = 'h5132;
    'h1476: romdata_int = 'h5c00;
    'h1477: romdata_int = 'h6280;
    'h1478: romdata_int = 'h78fd;
    'h1479: romdata_int = 'h7a41;
    'h147a: romdata_int = 'h8400;
    'h147b: romdata_int = 'ha937;
    'h147c: romdata_int = 'hac00;
    'h147d: romdata_int = 'hbe03;
    'h147e: romdata_int = 'hd400;
    'h147f: romdata_int = 'hd43d;
    'h1480: romdata_int = 'heaf2;
    'h1481: romdata_int = 'hfc00;
    'h1482: romdata_int = 'h100f0;
    'h1483: romdata_int = 'h10f09;
    'h1484: romdata_int = 'h11f37;
    'h1485: romdata_int = 'h12048;
    'h1486: romdata_int = 'h12400;
    'h1487: romdata_int = 'h5814; // Line descriptor for 8_9
    'h1488: romdata_int = 'h42e;
    'h1489: romdata_int = 'ha60;
    'h148a: romdata_int = 'he00;
    'h148b: romdata_int = 'h1328;
    'h148c: romdata_int = 'h2e9f;
    'h148d: romdata_int = 'h2f2d;
    'h148e: romdata_int = 'h3600;
    'h148f: romdata_int = 'h5e00;
    'h1490: romdata_int = 'h6c2b;
    'h1491: romdata_int = 'h76b0;
    'h1492: romdata_int = 'h814c;
    'h1493: romdata_int = 'h8600;
    'h1494: romdata_int = 'h8c32;
    'h1495: romdata_int = 'had56;
    'h1496: romdata_int = 'hae00;
    'h1497: romdata_int = 'hb069;
    'h1498: romdata_int = 'hd600;
    'h1499: romdata_int = 'he31d;
    'h149a: romdata_int = 'hef64;
    'h149b: romdata_int = 'hfe00;
    'h149c: romdata_int = 'hfeaa;
    'h149d: romdata_int = 'h1074b;
    'h149e: romdata_int = 'h11b49;
    'h149f: romdata_int = 'h122c3;
    'h14a0: romdata_int = 'h12600;
    'h14a1: romdata_int = 'h5814; // Line descriptor for 8_9
    'h14a2: romdata_int = 'h8e;
    'h14a3: romdata_int = 'h30b;
    'h14a4: romdata_int = 'h1000;
    'h14a5: romdata_int = 'h1079;
    'h14a6: romdata_int = 'h3800;
    'h14a7: romdata_int = 'h3a4f;
    'h14a8: romdata_int = 'h4ec5;
    'h14a9: romdata_int = 'h6000;
    'h14aa: romdata_int = 'h6661;
    'h14ab: romdata_int = 'h6946;
    'h14ac: romdata_int = 'h786b;
    'h14ad: romdata_int = 'h8800;
    'h14ae: romdata_int = 'h8cf6;
    'h14af: romdata_int = 'ha497;
    'h14b0: romdata_int = 'hb000;
    'h14b1: romdata_int = 'hb53f;
    'h14b2: romdata_int = 'hce3d;
    'h14b3: romdata_int = 'hd6e3;
    'h14b4: romdata_int = 'hd800;
    'h14b5: romdata_int = 'h10000;
    'h14b6: romdata_int = 'h1050b;
    'h14b7: romdata_int = 'h10afe;
    'h14b8: romdata_int = 'h12800;
    'h14b9: romdata_int = 'h12e5b;
    'h14ba: romdata_int = 'h13d1e;
    'h14bb: romdata_int = 'h5814; // Line descriptor for 8_9
    'h14bc: romdata_int = 'hd3b;
    'h14bd: romdata_int = 'h1200;
    'h14be: romdata_int = 'h1ab0;
    'h14bf: romdata_int = 'h1ce5;
    'h14c0: romdata_int = 'h3a00;
    'h14c1: romdata_int = 'h4262;
    'h14c2: romdata_int = 'h42c1;
    'h14c3: romdata_int = 'h525f;
    'h14c4: romdata_int = 'h6200;
    'h14c5: romdata_int = 'h643e;
    'h14c6: romdata_int = 'h8a00;
    'h14c7: romdata_int = 'h908f;
    'h14c8: romdata_int = 'h9d45;
    'h14c9: romdata_int = 'ha0a8;
    'h14ca: romdata_int = 'hb052;
    'h14cb: romdata_int = 'hb200;
    'h14cc: romdata_int = 'hda00;
    'h14cd: romdata_int = 'he8e4;
    'h14ce: romdata_int = 'he93e;
    'h14cf: romdata_int = 'hfca6;
    'h14d0: romdata_int = 'h10200;
    'h14d1: romdata_int = 'h10cc2;
    'h14d2: romdata_int = 'h128d5;
    'h14d3: romdata_int = 'h12a00;
    'h14d4: romdata_int = 'h13685;
    'h14d5: romdata_int = 'h5814; // Line descriptor for 8_9
    'h14d6: romdata_int = 'h404;
    'h14d7: romdata_int = 'he99;
    'h14d8: romdata_int = 'h1400;
    'h14d9: romdata_int = 'h1461;
    'h14da: romdata_int = 'h2c06;
    'h14db: romdata_int = 'h328f;
    'h14dc: romdata_int = 'h3c00;
    'h14dd: romdata_int = 'h542a;
    'h14de: romdata_int = 'h62ab;
    'h14df: romdata_int = 'h6400;
    'h14e0: romdata_int = 'h88c4;
    'h14e1: romdata_int = 'h8c00;
    'h14e2: romdata_int = 'h96dc;
    'h14e3: romdata_int = 'hb400;
    'h14e4: romdata_int = 'hbb60;
    'h14e5: romdata_int = 'hc094;
    'h14e6: romdata_int = 'hc830;
    'h14e7: romdata_int = 'hccf3;
    'h14e8: romdata_int = 'hdc00;
    'h14e9: romdata_int = 'hf487;
    'h14ea: romdata_int = 'hfa05;
    'h14eb: romdata_int = 'h10400;
    'h14ec: romdata_int = 'h12c00;
    'h14ed: romdata_int = 'h12e12;
    'h14ee: romdata_int = 'h1354e;
    'h14ef: romdata_int = 'h5814; // Line descriptor for 8_9
    'h14f0: romdata_int = 'h1600;
    'h14f1: romdata_int = 'h16ae;
    'h14f2: romdata_int = 'h203b;
    'h14f3: romdata_int = 'h2553;
    'h14f4: romdata_int = 'h3441;
    'h14f5: romdata_int = 'h3e00;
    'h14f6: romdata_int = 'h44b2;
    'h14f7: romdata_int = 'h5b06;
    'h14f8: romdata_int = 'h6040;
    'h14f9: romdata_int = 'h6600;
    'h14fa: romdata_int = 'h7c2b;
    'h14fb: romdata_int = 'h8a0a;
    'h14fc: romdata_int = 'h8e00;
    'h14fd: romdata_int = 'ha097;
    'h14fe: romdata_int = 'hb600;
    'h14ff: romdata_int = 'hbed8;
    'h1500: romdata_int = 'hd759;
    'h1501: romdata_int = 'hde00;
    'h1502: romdata_int = 'he111;
    'h1503: romdata_int = 'hf061;
    'h1504: romdata_int = 'h10600;
    'h1505: romdata_int = 'h11745;
    'h1506: romdata_int = 'h11c37;
    'h1507: romdata_int = 'h12e00;
    'h1508: romdata_int = 'h13b02;
    'h1509: romdata_int = 'h5814; // Line descriptor for 8_9
    'h150a: romdata_int = 'h2ae;
    'h150b: romdata_int = 'h83a;
    'h150c: romdata_int = 'h1800;
    'h150d: romdata_int = 'h1c6a;
    'h150e: romdata_int = 'h4000;
    'h150f: romdata_int = 'h4158;
    'h1510: romdata_int = 'h46e7;
    'h1511: romdata_int = 'h5c08;
    'h1512: romdata_int = 'h5c65;
    'h1513: romdata_int = 'h6800;
    'h1514: romdata_int = 'h84f6;
    'h1515: romdata_int = 'h9000;
    'h1516: romdata_int = 'h9250;
    'h1517: romdata_int = 'hae60;
    'h1518: romdata_int = 'hb800;
    'h1519: romdata_int = 'hc2e8;
    'h151a: romdata_int = 'hc880;
    'h151b: romdata_int = 'he000;
    'h151c: romdata_int = 'hed62;
    'h151d: romdata_int = 'h10800;
    'h151e: romdata_int = 'h10ad2;
    'h151f: romdata_int = 'h11627;
    'h1520: romdata_int = 'h12d3e;
    'h1521: romdata_int = 'h13000;
    'h1522: romdata_int = 'h13b2a;
    'h1523: romdata_int = 'h5814; // Line descriptor for 8_9
    'h1524: romdata_int = 'h101e;
    'h1525: romdata_int = 'h14d5;
    'h1526: romdata_int = 'h16e6;
    'h1527: romdata_int = 'h1a00;
    'h1528: romdata_int = 'h387d;
    'h1529: romdata_int = 'h4200;
    'h152a: romdata_int = 'h4a30;
    'h152b: romdata_int = 'h521c;
    'h152c: romdata_int = 'h6a00;
    'h152d: romdata_int = 'h6cba;
    'h152e: romdata_int = 'h9200;
    'h152f: romdata_int = 'h9232;
    'h1530: romdata_int = 'h942f;
    'h1531: romdata_int = 'haedd;
    'h1532: romdata_int = 'hba00;
    'h1533: romdata_int = 'hbcb4;
    'h1534: romdata_int = 'hcf59;
    'h1535: romdata_int = 'he0bd;
    'h1536: romdata_int = 'he200;
    'h1537: romdata_int = 'hf638;
    'h1538: romdata_int = 'h108fd;
    'h1539: romdata_int = 'h10a00;
    'h153a: romdata_int = 'h1248f;
    'h153b: romdata_int = 'h12656;
    'h153c: romdata_int = 'h13200;
    'h153d: romdata_int = 'h5814; // Line descriptor for 8_9
    'h153e: romdata_int = 'hcb9;
    'h153f: romdata_int = 'hf65;
    'h1540: romdata_int = 'h1c00;
    'h1541: romdata_int = 'h252c;
    'h1542: romdata_int = 'h3e66;
    'h1543: romdata_int = 'h4400;
    'h1544: romdata_int = 'h4ebd;
    'h1545: romdata_int = 'h54c9;
    'h1546: romdata_int = 'h6c00;
    'h1547: romdata_int = 'h6e44;
    'h1548: romdata_int = 'h8115;
    'h1549: romdata_int = 'h8a9a;
    'h154a: romdata_int = 'h9400;
    'h154b: romdata_int = 'haa36;
    'h154c: romdata_int = 'hb8b8;
    'h154d: romdata_int = 'hbc00;
    'h154e: romdata_int = 'hdc17;
    'h154f: romdata_int = 'hde6b;
    'h1550: romdata_int = 'he400;
    'h1551: romdata_int = 'hf8b8;
    'h1552: romdata_int = 'h1020a;
    'h1553: romdata_int = 'h10c00;
    'h1554: romdata_int = 'h118c4;
    'h1555: romdata_int = 'h13267;
    'h1556: romdata_int = 'h13400;
    'h1557: romdata_int = 'h5814; // Line descriptor for 8_9
    'h1558: romdata_int = 'h137;
    'h1559: romdata_int = 'hc7c;
    'h155a: romdata_int = 'h1cc9;
    'h155b: romdata_int = 'h1e00;
    'h155c: romdata_int = 'h3c1a;
    'h155d: romdata_int = 'h4600;
    'h155e: romdata_int = 'h48a0;
    'h155f: romdata_int = 'h5e5d;
    'h1560: romdata_int = 'h5e7b;
    'h1561: romdata_int = 'h6e00;
    'h1562: romdata_int = 'h8e3d;
    'h1563: romdata_int = 'h9600;
    'h1564: romdata_int = 'h96e3;
    'h1565: romdata_int = 'ha94c;
    'h1566: romdata_int = 'haaf4;
    'h1567: romdata_int = 'hbe00;
    'h1568: romdata_int = 'hd413;
    'h1569: romdata_int = 'he24f;
    'h156a: romdata_int = 'he600;
    'h156b: romdata_int = 'hfa43;
    'h156c: romdata_int = 'h10e00;
    'h156d: romdata_int = 'h1143b;
    'h156e: romdata_int = 'h12718;
    'h156f: romdata_int = 'h130ea;
    'h1570: romdata_int = 'h13600;
    'h1571: romdata_int = 'h5814; // Line descriptor for 8_9
    'h1572: romdata_int = 'h6e1;
    'h1573: romdata_int = 'h1455;
    'h1574: romdata_int = 'h2000;
    'h1575: romdata_int = 'h2549;
    'h1576: romdata_int = 'h2901;
    'h1577: romdata_int = 'h2ad9;
    'h1578: romdata_int = 'h4800;
    'h1579: romdata_int = 'h509f;
    'h157a: romdata_int = 'h6ab4;
    'h157b: romdata_int = 'h7000;
    'h157c: romdata_int = 'h86ed;
    'h157d: romdata_int = 'h873d;
    'h157e: romdata_int = 'h9800;
    'h157f: romdata_int = 'hc000;
    'h1580: romdata_int = 'hc059;
    'h1581: romdata_int = 'hc71e;
    'h1582: romdata_int = 'hd291;
    'h1583: romdata_int = 'he800;
    'h1584: romdata_int = 'hea2c;
    'h1585: romdata_int = 'hfd50;
    'h1586: romdata_int = 'h102d2;
    'h1587: romdata_int = 'h11000;
    'h1588: romdata_int = 'h11d49;
    'h1589: romdata_int = 'h13800;
    'h158a: romdata_int = 'h13e54;
    'h158b: romdata_int = 'h5814; // Line descriptor for 8_9
    'h158c: romdata_int = 'h489;
    'h158d: romdata_int = 'h8a1;
    'h158e: romdata_int = 'h1f50;
    'h158f: romdata_int = 'h2200;
    'h1590: romdata_int = 'h394a;
    'h1591: romdata_int = 'h4a00;
    'h1592: romdata_int = 'h4a9b;
    'h1593: romdata_int = 'h6018;
    'h1594: romdata_int = 'h7200;
    'h1595: romdata_int = 'h72c3;
    'h1596: romdata_int = 'h8323;
    'h1597: romdata_int = 'h9a00;
    'h1598: romdata_int = 'h9c78;
    'h1599: romdata_int = 'ha2b1;
    'h159a: romdata_int = 'hc200;
    'h159b: romdata_int = 'hc4ee;
    'h159c: romdata_int = 'hcce5;
    'h159d: romdata_int = 'hd033;
    'h159e: romdata_int = 'hea00;
    'h159f: romdata_int = 'hf29b;
    'h15a0: romdata_int = 'hf820;
    'h15a1: romdata_int = 'h11200;
    'h15a2: romdata_int = 'h11e48;
    'h15a3: romdata_int = 'h13644;
    'h15a4: romdata_int = 'h13a00;
    'h15a5: romdata_int = 'h5814; // Line descriptor for 8_9
    'h15a6: romdata_int = 'h212b;
    'h15a7: romdata_int = 'h2400;
    'h15a8: romdata_int = 'h2688;
    'h15a9: romdata_int = 'h2727;
    'h15aa: romdata_int = 'h314f;
    'h15ab: romdata_int = 'h4c00;
    'h15ac: romdata_int = 'h4d35;
    'h15ad: romdata_int = 'h70ea;
    'h15ae: romdata_int = 'h7400;
    'h15af: romdata_int = 'h74ca;
    'h15b0: romdata_int = 'h8814;
    'h15b1: romdata_int = 'h9b20;
    'h15b2: romdata_int = 'h9c00;
    'h15b3: romdata_int = 'ha6a2;
    'h15b4: romdata_int = 'hc2a0;
    'h15b5: romdata_int = 'hc400;
    'h15b6: romdata_int = 'hd8e6;
    'h15b7: romdata_int = 'hdf15;
    'h15b8: romdata_int = 'hec00;
    'h15b9: romdata_int = 'hf13d;
    'h15ba: romdata_int = 'h10e17;
    'h15bb: romdata_int = 'h11400;
    'h15bc: romdata_int = 'h1188a;
    'h15bd: romdata_int = 'h11aa1;
    'h15be: romdata_int = 'h13c00;
    'h15bf: romdata_int = 'h7814; // Line descriptor for 8_9
    'h15c0: romdata_int = 'h6ec;
    'h15c1: romdata_int = 'h1734;
    'h15c2: romdata_int = 'h1e4e;
    'h15c3: romdata_int = 'h2600;
    'h15c4: romdata_int = 'h3025;
    'h15c5: romdata_int = 'h3633;
    'h15c6: romdata_int = 'h4e00;
    'h15c7: romdata_int = 'h6890;
    'h15c8: romdata_int = 'h745c;
    'h15c9: romdata_int = 'h7600;
    'h15ca: romdata_int = 'h7c73;
    'h15cb: romdata_int = 'h8210;
    'h15cc: romdata_int = 'h9e00;
    'h15cd: romdata_int = 'hb269;
    'h15ce: romdata_int = 'hc600;
    'h15cf: romdata_int = 'hc645;
    'h15d0: romdata_int = 'hcb49;
    'h15d1: romdata_int = 'hd0cf;
    'h15d2: romdata_int = 'hee00;
    'h15d3: romdata_int = 'h10518;
    'h15d4: romdata_int = 'h1151c;
    'h15d5: romdata_int = 'h11600;
    'h15d6: romdata_int = 'h12555;
    'h15d7: romdata_int = 'h13e00;
    'h15d8: romdata_int = 'h13e48;
    'h15d9: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h15da: romdata_int = 'h0;
    'h15db: romdata_int = 'h322;
    'h15dc: romdata_int = 'h172c;
    'h15dd: romdata_int = 'h1ac4;
    'h15de: romdata_int = 'h2400;
    'h15df: romdata_int = 'h3538;
    'h15e0: romdata_int = 'h4679;
    'h15e1: romdata_int = 'h4800;
    'h15e2: romdata_int = 'h4ad0;
    'h15e3: romdata_int = 'h6a7e;
    'h15e4: romdata_int = 'h6c00;
    'h15e5: romdata_int = 'h7272;
    'h15e6: romdata_int = 'h8123;
    'h15e7: romdata_int = 'h9000;
    'h15e8: romdata_int = 'ha84a;
    'h15e9: romdata_int = 'hac67;
    'h15ea: romdata_int = 'hb400;
    'h15eb: romdata_int = 'hb608;
    'h15ec: romdata_int = 'hc2ed;
    'h15ed: romdata_int = 'hd800;
    'h15ee: romdata_int = 'he15c;
    'h15ef: romdata_int = 'hf8d8;
    'h15f0: romdata_int = 'hfc00;
    'h15f1: romdata_int = 'hfc5e;
    'h15f2: romdata_int = 'h1063a;
    'h15f3: romdata_int = 'h12000;
    'h15f4: romdata_int = 'h13241;
    'h15f5: romdata_int = 'h13440;
    'h15f6: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h15f7: romdata_int = 'h200;
    'h15f8: romdata_int = 'h75c;
    'h15f9: romdata_int = 'hebc;
    'h15fa: romdata_int = 'h1928;
    'h15fb: romdata_int = 'h2600;
    'h15fc: romdata_int = 'h3d05;
    'h15fd: romdata_int = 'h3f48;
    'h15fe: romdata_int = 'h4a00;
    'h15ff: romdata_int = 'h5850;
    'h1600: romdata_int = 'h5919;
    'h1601: romdata_int = 'h6e00;
    'h1602: romdata_int = 'h70eb;
    'h1603: romdata_int = 'h7cad;
    'h1604: romdata_int = 'h9200;
    'h1605: romdata_int = 'h961e;
    'h1606: romdata_int = 'haec8;
    'h1607: romdata_int = 'hb600;
    'h1608: romdata_int = 'hbc67;
    'h1609: romdata_int = 'hc8d6;
    'h160a: romdata_int = 'hda00;
    'h160b: romdata_int = 'hed28;
    'h160c: romdata_int = 'hee24;
    'h160d: romdata_int = 'hfe00;
    'h160e: romdata_int = 'h11824;
    'h160f: romdata_int = 'h11eea;
    'h1610: romdata_int = 'h12141;
    'h1611: romdata_int = 'h12200;
    'h1612: romdata_int = 'h13d2c;
    'h1613: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h1614: romdata_int = 'ha1;
    'h1615: romdata_int = 'h400;
    'h1616: romdata_int = 'h100d;
    'h1617: romdata_int = 'h204a;
    'h1618: romdata_int = 'h2800;
    'h1619: romdata_int = 'h3675;
    'h161a: romdata_int = 'h44c1;
    'h161b: romdata_int = 'h4831;
    'h161c: romdata_int = 'h4c00;
    'h161d: romdata_int = 'h50bd;
    'h161e: romdata_int = 'h7000;
    'h161f: romdata_int = 'h74ee;
    'h1620: romdata_int = 'h7c35;
    'h1621: romdata_int = 'h9400;
    'h1622: romdata_int = 'h9ee5;
    'h1623: romdata_int = 'ha4f3;
    'h1624: romdata_int = 'hb800;
    'h1625: romdata_int = 'hc470;
    'h1626: romdata_int = 'hc8ce;
    'h1627: romdata_int = 'hdb21;
    'h1628: romdata_int = 'hdc00;
    'h1629: romdata_int = 'hf932;
    'h162a: romdata_int = 'h10000;
    'h162b: romdata_int = 'h11304;
    'h162c: romdata_int = 'h11e50;
    'h162d: romdata_int = 'h12400;
    'h162e: romdata_int = 'h12454;
    'h162f: romdata_int = 'h13f1a;
    'h1630: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h1631: romdata_int = 'h600;
    'h1632: romdata_int = 'hab8;
    'h1633: romdata_int = 'h1843;
    'h1634: romdata_int = 'h2077;
    'h1635: romdata_int = 'h28bd;
    'h1636: romdata_int = 'h2a00;
    'h1637: romdata_int = 'h2e5f;
    'h1638: romdata_int = 'h4e00;
    'h1639: romdata_int = 'h4ebe;
    'h163a: romdata_int = 'h6825;
    'h163b: romdata_int = 'h7200;
    'h163c: romdata_int = 'h8ab3;
    'h163d: romdata_int = 'h8e32;
    'h163e: romdata_int = 'h9600;
    'h163f: romdata_int = 'h9c1d;
    'h1640: romdata_int = 'h9e3c;
    'h1641: romdata_int = 'hba00;
    'h1642: romdata_int = 'hd246;
    'h1643: romdata_int = 'hd503;
    'h1644: romdata_int = 'hd8b0;
    'h1645: romdata_int = 'hdd35;
    'h1646: romdata_int = 'hde00;
    'h1647: romdata_int = 'h10200;
    'h1648: romdata_int = 'h10eca;
    'h1649: romdata_int = 'h114a9;
    'h164a: romdata_int = 'h1247b;
    'h164b: romdata_int = 'h12600;
    'h164c: romdata_int = 'h1304b;
    'h164d: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h164e: romdata_int = 'h800;
    'h164f: romdata_int = 'h939;
    'h1650: romdata_int = 'ha79;
    'h1651: romdata_int = 'h1c52;
    'h1652: romdata_int = 'h2c00;
    'h1653: romdata_int = 'h2c4b;
    'h1654: romdata_int = 'h309f;
    'h1655: romdata_int = 'h5000;
    'h1656: romdata_int = 'h5a21;
    'h1657: romdata_int = 'h6680;
    'h1658: romdata_int = 'h7400;
    'h1659: romdata_int = 'h7a41;
    'h165a: romdata_int = 'h88f6;
    'h165b: romdata_int = 'h9800;
    'h165c: romdata_int = 'h9aa1;
    'h165d: romdata_int = 'ha081;
    'h165e: romdata_int = 'hb462;
    'h165f: romdata_int = 'hb4b4;
    'h1660: romdata_int = 'hbc00;
    'h1661: romdata_int = 'he000;
    'h1662: romdata_int = 'he4b4;
    'h1663: romdata_int = 'he6df;
    'h1664: romdata_int = 'hfd44;
    'h1665: romdata_int = 'h10400;
    'h1666: romdata_int = 'h10cc2;
    'h1667: romdata_int = 'h12800;
    'h1668: romdata_int = 'h13115;
    'h1669: romdata_int = 'h1372a;
    'h166a: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h166b: romdata_int = 'ha00;
    'h166c: romdata_int = 'h1091;
    'h166d: romdata_int = 'h16a4;
    'h166e: romdata_int = 'h20e7;
    'h166f: romdata_int = 'h252c;
    'h1670: romdata_int = 'h2e00;
    'h1671: romdata_int = 'h40ee;
    'h1672: romdata_int = 'h5200;
    'h1673: romdata_int = 'h5c1a;
    'h1674: romdata_int = 'h5d2c;
    'h1675: romdata_int = 'h7600;
    'h1676: romdata_int = 'h7733;
    'h1677: romdata_int = 'h7a07;
    'h1678: romdata_int = 'h94f2;
    'h1679: romdata_int = 'h94f6;
    'h167a: romdata_int = 'h9a00;
    'h167b: romdata_int = 'hb858;
    'h167c: romdata_int = 'hbe00;
    'h167d: romdata_int = 'hd210;
    'h167e: romdata_int = 'he200;
    'h167f: romdata_int = 'hf2d3;
    'h1680: romdata_int = 'hf4ad;
    'h1681: romdata_int = 'h10600;
    'h1682: romdata_int = 'h1095f;
    'h1683: romdata_int = 'h10b37;
    'h1684: romdata_int = 'h12a00;
    'h1685: romdata_int = 'h12a54;
    'h1686: romdata_int = 'h13e95;
    'h1687: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h1688: romdata_int = 'h42e;
    'h1689: romdata_int = 'ha60;
    'h168a: romdata_int = 'hc00;
    'h168b: romdata_int = 'h1128;
    'h168c: romdata_int = 'h26a6;
    'h168d: romdata_int = 'h2b34;
    'h168e: romdata_int = 'h3000;
    'h168f: romdata_int = 'h50c5;
    'h1690: romdata_int = 'h5400;
    'h1691: romdata_int = 'h683e;
    'h1692: romdata_int = 'h7800;
    'h1693: romdata_int = 'h78fd;
    'h1694: romdata_int = 'h8832;
    'h1695: romdata_int = 'h9c00;
    'h1696: romdata_int = 'h9c97;
    'h1697: romdata_int = 'haf3f;
    'h1698: romdata_int = 'hbb1e;
    'h1699: romdata_int = 'hbe96;
    'h169a: romdata_int = 'hc000;
    'h169b: romdata_int = 'he291;
    'h169c: romdata_int = 'he400;
    'h169d: romdata_int = 'hf317;
    'h169e: romdata_int = 'h10800;
    'h169f: romdata_int = 'h10ec3;
    'h16a0: romdata_int = 'h11691;
    'h16a1: romdata_int = 'h128d6;
    'h16a2: romdata_int = 'h12c00;
    'h16a3: romdata_int = 'h12f25;
    'h16a4: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h16a5: romdata_int = 'h8e;
    'h16a6: romdata_int = 'h30b;
    'h16a7: romdata_int = 'he00;
    'h16a8: romdata_int = 'he79;
    'h16a9: romdata_int = 'h312d;
    'h16aa: romdata_int = 'h3200;
    'h16ab: romdata_int = 'h3911;
    'h16ac: romdata_int = 'h48e7;
    'h16ad: romdata_int = 'h5332;
    'h16ae: romdata_int = 'h5600;
    'h16af: romdata_int = 'h7044;
    'h16b0: romdata_int = 'h74c3;
    'h16b1: romdata_int = 'h7a00;
    'h16b2: romdata_int = 'h9e00;
    'h16b3: romdata_int = 'ha337;
    'h16b4: romdata_int = 'ha956;
    'h16b5: romdata_int = 'hb677;
    'h16b6: romdata_int = 'hb8ee;
    'h16b7: romdata_int = 'hc200;
    'h16b8: romdata_int = 'he600;
    'h16b9: romdata_int = 'he87d;
    'h16ba: romdata_int = 'he8aa;
    'h16bb: romdata_int = 'h10a00;
    'h16bc: romdata_int = 'h10c48;
    'h16bd: romdata_int = 'h1107f;
    'h16be: romdata_int = 'h1291e;
    'h16bf: romdata_int = 'h12e00;
    'h16c0: romdata_int = 'h1384e;
    'h16c1: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h16c2: romdata_int = 'hd3b;
    'h16c3: romdata_int = 'h1000;
    'h16c4: romdata_int = 'h16f3;
    'h16c5: romdata_int = 'h220e;
    'h16c6: romdata_int = 'h3400;
    'h16c7: romdata_int = 'h348f;
    'h16c8: romdata_int = 'h3c4f;
    'h16c9: romdata_int = 'h5800;
    'h16ca: romdata_int = 'h5f06;
    'h16cb: romdata_int = 'h5f21;
    'h16cc: romdata_int = 'h6e2b;
    'h16cd: romdata_int = 'h7c00;
    'h16ce: romdata_int = 'h7e3c;
    'h16cf: romdata_int = 'ha000;
    'h16d0: romdata_int = 'hb0b5;
    'h16d1: romdata_int = 'hb150;
    'h16d2: romdata_int = 'hc400;
    'h16d3: romdata_int = 'hcd55;
    'h16d4: romdata_int = 'hd762;
    'h16d5: romdata_int = 'hda75;
    'h16d6: romdata_int = 'he800;
    'h16d7: romdata_int = 'hec42;
    'h16d8: romdata_int = 'h10652;
    'h16d9: romdata_int = 'h10c00;
    'h16da: romdata_int = 'h11b5a;
    'h16db: romdata_int = 'h12caf;
    'h16dc: romdata_int = 'h13000;
    'h16dd: romdata_int = 'h142bc;
    'h16de: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h16df: romdata_int = 'h404;
    'h16e0: romdata_int = 'h1200;
    'h16e1: romdata_int = 'h1261;
    'h16e2: romdata_int = 'h1ed5;
    'h16e3: romdata_int = 'h2e06;
    'h16e4: romdata_int = 'h3600;
    'h16e5: romdata_int = 'h3641;
    'h16e6: romdata_int = 'h545f;
    'h16e7: romdata_int = 'h562a;
    'h16e8: romdata_int = 'h5a00;
    'h16e9: romdata_int = 'h786b;
    'h16ea: romdata_int = 'h7e00;
    'h16eb: romdata_int = 'h8c8f;
    'h16ec: romdata_int = 'h902f;
    'h16ed: romdata_int = 'ha14d;
    'h16ee: romdata_int = 'ha200;
    'h16ef: romdata_int = 'hc226;
    'h16f0: romdata_int = 'hc600;
    'h16f1: romdata_int = 'hd54a;
    'h16f2: romdata_int = 'hea00;
    'h16f3: romdata_int = 'hf0fe;
    'h16f4: romdata_int = 'hf709;
    'h16f5: romdata_int = 'h10156;
    'h16f6: romdata_int = 'h10e00;
    'h16f7: romdata_int = 'h118b5;
    'h16f8: romdata_int = 'h12285;
    'h16f9: romdata_int = 'h13200;
    'h16fa: romdata_int = 'h14061;
    'h16fb: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h16fc: romdata_int = 'h1400;
    'h16fd: romdata_int = 'h14ae;
    'h16fe: romdata_int = 'h1c3b;
    'h16ff: romdata_int = 'h2283;
    'h1700: romdata_int = 'h3800;
    'h1701: romdata_int = 'h4066;
    'h1702: romdata_int = 'h432a;
    'h1703: romdata_int = 'h4c30;
    'h1704: romdata_int = 'h5c00;
    'h1705: romdata_int = 'h66ab;
    'h1706: romdata_int = 'h6d46;
    'h1707: romdata_int = 'h8000;
    'h1708: romdata_int = 'h869a;
    'h1709: romdata_int = 'h92dc;
    'h170a: romdata_int = 'ha400;
    'h170b: romdata_int = 'hb2b8;
    'h170c: romdata_int = 'hba45;
    'h170d: romdata_int = 'hc800;
    'h170e: romdata_int = 'hd11d;
    'h170f: romdata_int = 'hd904;
    'h1710: romdata_int = 'he438;
    'h1711: romdata_int = 'hec00;
    'h1712: romdata_int = 'h108e0;
    'h1713: romdata_int = 'h11000;
    'h1714: romdata_int = 'h1169c;
    'h1715: romdata_int = 'h13400;
    'h1716: romdata_int = 'h134f2;
    'h1717: romdata_int = 'h14011;
    'h1718: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h1719: romdata_int = 'h2ae;
    'h171a: romdata_int = 'h83a;
    'h171b: romdata_int = 'h1600;
    'h171c: romdata_int = 'h18b0;
    'h171d: romdata_int = 'h3a00;
    'h171e: romdata_int = 'h3a7d;
    'h171f: romdata_int = 'h4462;
    'h1720: romdata_int = 'h4c9b;
    'h1721: romdata_int = 'h5e00;
    'h1722: romdata_int = 'h6008;
    'h1723: romdata_int = 'h6eba;
    'h1724: romdata_int = 'h8200;
    'h1725: romdata_int = 'h860a;
    'h1726: romdata_int = 'h90f8;
    'h1727: romdata_int = 'h92e3;
    'h1728: romdata_int = 'ha600;
    'h1729: romdata_int = 'hca00;
    'h172a: romdata_int = 'hcb1c;
    'h172b: romdata_int = 'hccb8;
    'h172c: romdata_int = 'hde61;
    'h172d: romdata_int = 'hee00;
    'h172e: romdata_int = 'hf0d2;
    'h172f: romdata_int = 'h1047b;
    'h1730: romdata_int = 'h11200;
    'h1731: romdata_int = 'h112d5;
    'h1732: romdata_int = 'h12737;
    'h1733: romdata_int = 'h13600;
    'h1734: romdata_int = 'h1426e;
    'h1735: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h1736: romdata_int = 'hcb9;
    'h1737: romdata_int = 'he1e;
    'h1738: romdata_int = 'h12d5;
    'h1739: romdata_int = 'h1800;
    'h173a: romdata_int = 'h3c00;
    'h173b: romdata_int = 'h3e1a;
    'h173c: romdata_int = 'h46b2;
    'h173d: romdata_int = 'h541c;
    'h173e: romdata_int = 'h6000;
    'h173f: romdata_int = 'h6440;
    'h1740: romdata_int = 'h80f6;
    'h1741: romdata_int = 'h8400;
    'h1742: romdata_int = 'h84c4;
    'h1743: romdata_int = 'h983f;
    'h1744: romdata_int = 'ha636;
    'h1745: romdata_int = 'ha800;
    'h1746: romdata_int = 'hc0ba;
    'h1747: romdata_int = 'hcc00;
    'h1748: romdata_int = 'hd6fc;
    'h1749: romdata_int = 'hdd62;
    'h174a: romdata_int = 'heed9;
    'h174b: romdata_int = 'hf000;
    'h174c: romdata_int = 'h102c4;
    'h174d: romdata_int = 'h10560;
    'h174e: romdata_int = 'h11400;
    'h174f: romdata_int = 'h12058;
    'h1750: romdata_int = 'h13800;
    'h1751: romdata_int = 'h13c55;
    'h1752: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h1753: romdata_int = 'h137;
    'h1754: romdata_int = 'h1a00;
    'h1755: romdata_int = 'h1e62;
    'h1756: romdata_int = 'h1ef2;
    'h1757: romdata_int = 'h285c;
    'h1758: romdata_int = 'h3b4a;
    'h1759: romdata_int = 'h3e00;
    'h175a: romdata_int = 'h56c9;
    'h175b: romdata_int = 'h5b38;
    'h175c: romdata_int = 'h6200;
    'h175d: romdata_int = 'h72ea;
    'h175e: romdata_int = 'h8600;
    'h175f: romdata_int = 'h8a3d;
    'h1760: romdata_int = 'ha457;
    'h1761: romdata_int = 'haa00;
    'h1762: romdata_int = 'hab29;
    'h1763: romdata_int = 'hca33;
    'h1764: romdata_int = 'hce00;
    'h1765: romdata_int = 'hce6b;
    'h1766: romdata_int = 'heaaa;
    'h1767: romdata_int = 'hf200;
    'h1768: romdata_int = 'hfaf3;
    'h1769: romdata_int = 'h1111e;
    'h176a: romdata_int = 'h11423;
    'h176b: romdata_int = 'h11600;
    'h176c: romdata_int = 'h12244;
    'h176d: romdata_int = 'h13a00;
    'h176e: romdata_int = 'h13b39;
    'h176f: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h1770: romdata_int = 'h6e1;
    'h1771: romdata_int = 'hc7c;
    'h1772: romdata_int = 'h14e6;
    'h1773: romdata_int = 'h1c00;
    'h1774: romdata_int = 'h26f2;
    'h1775: romdata_int = 'h2b01;
    'h1776: romdata_int = 'h4000;
    'h1777: romdata_int = 'h529f;
    'h1778: romdata_int = 'h6065;
    'h1779: romdata_int = 'h6400;
    'h177a: romdata_int = 'h82ed;
    'h177b: romdata_int = 'h8800;
    'h177c: romdata_int = 'h8d5d;
    'h177d: romdata_int = 'h9720;
    'h177e: romdata_int = 'ha34c;
    'h177f: romdata_int = 'hac00;
    'h1780: romdata_int = 'hbf0b;
    'h1781: romdata_int = 'hc629;
    'h1782: romdata_int = 'hd000;
    'h1783: romdata_int = 'he242;
    'h1784: romdata_int = 'hf400;
    'h1785: romdata_int = 'hf4c2;
    'h1786: romdata_int = 'hff1c;
    'h1787: romdata_int = 'h11800;
    'h1788: romdata_int = 'h11ca3;
    'h1789: romdata_int = 'h12627;
    'h178a: romdata_int = 'h13339;
    'h178b: romdata_int = 'h13c00;
    'h178c: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h178d: romdata_int = 'h489;
    'h178e: romdata_int = 'h1b50;
    'h178f: romdata_int = 'h1e00;
    'h1790: romdata_int = 'h2318;
    'h1791: romdata_int = 'h2cd9;
    'h1792: romdata_int = 'h3833;
    'h1793: romdata_int = 'h4200;
    'h1794: romdata_int = 'h625d;
    'h1795: romdata_int = 'h627b;
    'h1796: romdata_int = 'h6600;
    'h1797: romdata_int = 'h7ead;
    'h1798: romdata_int = 'h8414;
    'h1799: romdata_int = 'h8a00;
    'h179a: romdata_int = 'ha6f4;
    'h179b: romdata_int = 'haadc;
    'h179c: romdata_int = 'hae00;
    'h179d: romdata_int = 'hc674;
    'h179e: romdata_int = 'hd04f;
    'h179f: romdata_int = 'hd200;
    'h17a0: romdata_int = 'he09b;
    'h17a1: romdata_int = 'he725;
    'h17a2: romdata_int = 'hf600;
    'h17a3: romdata_int = 'h1013d;
    'h17a4: romdata_int = 'h1028a;
    'h17a5: romdata_int = 'h11a00;
    'h17a6: romdata_int = 'h12e92;
    'h17a7: romdata_int = 'h136c5;
    'h17a8: romdata_int = 'h13e00;
    'h17a9: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h17aa: romdata_int = 'h8a1;
    'h17ab: romdata_int = 'h1255;
    'h17ac: romdata_int = 'h1d2b;
    'h17ad: romdata_int = 'h2000;
    'h17ae: romdata_int = 'h2553;
    'h17af: romdata_int = 'h4358;
    'h17b0: romdata_int = 'h4400;
    'h17b1: romdata_int = 'h4aa0;
    'h17b2: romdata_int = 'h6800;
    'h17b3: romdata_int = 'h6b3f;
    'h17b4: romdata_int = 'h76b0;
    'h17b5: romdata_int = 'h833d;
    'h17b6: romdata_int = 'h8c00;
    'h17b7: romdata_int = 'h98f5;
    'h17b8: romdata_int = 'h9ab1;
    'h17b9: romdata_int = 'hb000;
    'h17ba: romdata_int = 'hc4e6;
    'h17bb: romdata_int = 'hcf15;
    'h17bc: romdata_int = 'hd400;
    'h17bd: romdata_int = 'hdf3d;
    'h17be: romdata_int = 'hf800;
    'h17bf: romdata_int = 'hfae2;
    'h17c0: romdata_int = 'hfe3b;
    'h17c1: romdata_int = 'h11c00;
    'h17c2: romdata_int = 'h11c23;
    'h17c3: romdata_int = 'h12a48;
    'h17c4: romdata_int = 'h12c8d;
    'h17c5: romdata_int = 'h14000;
    'h17c6: romdata_int = 'h7b12; // Line descriptor for 9_10
    'h17c7: romdata_int = 'h6ec;
    'h17c8: romdata_int = 'h1534;
    'h17c9: romdata_int = 'h1a4e;
    'h17ca: romdata_int = 'h2200;
    'h17cb: romdata_int = 'h3225;
    'h17cc: romdata_int = 'h334f;
    'h17cd: romdata_int = 'h4600;
    'h17ce: romdata_int = 'h4f35;
    'h17cf: romdata_int = 'h6418;
    'h17d0: romdata_int = 'h6a00;
    'h17d1: romdata_int = 'h6c90;
    'h17d2: romdata_int = 'h8e00;
    'h17d3: romdata_int = 'h8e50;
    'h17d4: romdata_int = 'hac69;
    'h17d5: romdata_int = 'hb200;
    'h17d6: romdata_int = 'hb2e2;
    'h17d7: romdata_int = 'hbd49;
    'h17d8: romdata_int = 'hc051;
    'h17d9: romdata_int = 'hd600;
    'h17da: romdata_int = 'hea89;
    'h17db: romdata_int = 'hf617;
    'h17dc: romdata_int = 'hfa00;
    'h17dd: romdata_int = 'h10a48;
    'h17de: romdata_int = 'h11a20;
    'h17df: romdata_int = 'h11e00;
    'h17e0: romdata_int = 'h138c6;
    'h17e1: romdata_int = 'h13b02;
    'h17e2: romdata_int = 'h14200;
    'h17e3: romdata_int = 'h4124; // Line descriptor for 1_5s
    'h17e4: romdata_int = 'h667;
    'h17e5: romdata_int = 'h4;
    'h17e6: romdata_int = 'h124; // Line descriptor for 1_5s
    'h17e7: romdata_int = 'h6bd;
    'h17e8: romdata_int = 'ha5e;
    'h17e9: romdata_int = 'h124; // Line descriptor for 1_5s
    'h17ea: romdata_int = 'h261;
    'h17eb: romdata_int = 'h334;
    'h17ec: romdata_int = 'h124; // Line descriptor for 1_5s
    'h17ed: romdata_int = 'h4c9;
    'h17ee: romdata_int = 'he41;
    'h17ef: romdata_int = 'h124; // Line descriptor for 1_5s
    'h17f0: romdata_int = 'h2e;
    'h17f1: romdata_int = 'h89;
    'h17f2: romdata_int = 'h124; // Line descriptor for 1_5s
    'h17f3: romdata_int = 'h6a6;
    'h17f4: romdata_int = 'h2e0;
    'h17f5: romdata_int = 'h24; // Line descriptor for 1_5s
    'h17f6: romdata_int = 'h6f2;
    'h17f7: romdata_int = 'h4124; // Line descriptor for 1_5s
    'h17f8: romdata_int = 'h137;
    'h17f9: romdata_int = 'h26b;
    'h17fa: romdata_int = 'h124; // Line descriptor for 1_5s
    'h17fb: romdata_int = 'h4d5;
    'h17fc: romdata_int = 'h477;
    'h17fd: romdata_int = 'h124; // Line descriptor for 1_5s
    'h17fe: romdata_int = 'h92b;
    'h17ff: romdata_int = 'h108a;
    'h1800: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1801: romdata_int = 'h44a;
    'h1802: romdata_int = 'h52b;
    'h1803: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1804: romdata_int = 'hb0;
    'h1805: romdata_int = 'h255;
    'h1806: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1807: romdata_int = 'h688;
    'h1808: romdata_int = 'h1111;
    'h1809: romdata_int = 'h24; // Line descriptor for 1_5s
    'h180a: romdata_int = 'h464;
    'h180b: romdata_int = 'h24; // Line descriptor for 1_5s
    'h180c: romdata_int = 'h10b;
    'h180d: romdata_int = 'h4024; // Line descriptor for 1_5s
    'h180e: romdata_int = 'h86;
    'h180f: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1810: romdata_int = 'h8;
    'h1811: romdata_int = 'h2e6;
    'h1812: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1813: romdata_int = 'h536;
    'h1814: romdata_int = 'h31e;
    'h1815: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1816: romdata_int = 'hb2d;
    'h1817: romdata_int = 'h1161;
    'h1818: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1819: romdata_int = 'h855;
    'h181a: romdata_int = 'h2d5;
    'h181b: romdata_int = 'h24; // Line descriptor for 1_5s
    'h181c: romdata_int = 'h28a;
    'h181d: romdata_int = 'h124; // Line descriptor for 1_5s
    'h181e: romdata_int = 'h722;
    'h181f: romdata_int = 'h462;
    'h1820: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1821: romdata_int = 'hd4d;
    'h1822: romdata_int = 'h65c;
    'h1823: romdata_int = 'h4124; // Line descriptor for 1_5s
    'h1824: romdata_int = 'h9a;
    'h1825: romdata_int = 'ha9f;
    'h1826: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1827: romdata_int = 'h490;
    'h1828: romdata_int = 'h2a5;
    'h1829: romdata_int = 'h124; // Line descriptor for 1_5s
    'h182a: romdata_int = 'h554;
    'h182b: romdata_int = 'h749;
    'h182c: romdata_int = 'h24; // Line descriptor for 1_5s
    'h182d: romdata_int = 'h267;
    'h182e: romdata_int = 'h24; // Line descriptor for 1_5s
    'h182f: romdata_int = 'hd5;
    'h1830: romdata_int = 'h24; // Line descriptor for 1_5s
    'h1831: romdata_int = 'hc25;
    'h1832: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1833: romdata_int = 'h15c;
    'h1834: romdata_int = 'he75;
    'h1835: romdata_int = 'h24; // Line descriptor for 1_5s
    'h1836: romdata_int = 'h727;
    'h1837: romdata_int = 'h4124; // Line descriptor for 1_5s
    'h1838: romdata_int = 'h4b6;
    'h1839: romdata_int = 'hae;
    'h183a: romdata_int = 'h124; // Line descriptor for 1_5s
    'h183b: romdata_int = 'h8d9;
    'h183c: romdata_int = 'h734;
    'h183d: romdata_int = 'h124; // Line descriptor for 1_5s
    'h183e: romdata_int = 'heab;
    'h183f: romdata_int = 'h701;
    'h1840: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1841: romdata_int = 'h4f2;
    'h1842: romdata_int = 'hd52;
    'h1843: romdata_int = 'h2124; // Line descriptor for 1_5s
    'h1844: romdata_int = 'h328;
    'h1845: romdata_int = 'h648;
    'h1846: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1847: romdata_int = 'h48f;
    'h1848: romdata_int = 'h680;
    'h1849: romdata_int = 'h154b;
    'h184a: romdata_int = 'h421e; // Line descriptor for 1_3s
    'h184b: romdata_int = 'h91d;
    'h184c: romdata_int = 'h2c9;
    'h184d: romdata_int = 'h83d;
    'h184e: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h184f: romdata_int = 'h95d;
    'h1850: romdata_int = 'hcef;
    'h1851: romdata_int = 'h61;
    'h1852: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1853: romdata_int = 'h67b;
    'h1854: romdata_int = 'h12fc;
    'h1855: romdata_int = 'he0;
    'h1856: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1857: romdata_int = 'h425;
    'h1858: romdata_int = 'h1839;
    'h1859: romdata_int = 'h1c6f;
    'h185a: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h185b: romdata_int = 'ha32;
    'h185c: romdata_int = 'h277;
    'h185d: romdata_int = 'h6cf;
    'h185e: romdata_int = 'h421e; // Line descriptor for 1_3s
    'h185f: romdata_int = 'h2d5;
    'h1860: romdata_int = 'h6b;
    'h1861: romdata_int = 'h24a;
    'h1862: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1863: romdata_int = 'h552;
    'h1864: romdata_int = 'h65d;
    'h1865: romdata_int = 'h165a;
    'h1866: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1867: romdata_int = 'h32b;
    'h1868: romdata_int = 'hb03;
    'h1869: romdata_int = 'h1a81;
    'h186a: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h186b: romdata_int = 'h4ab;
    'h186c: romdata_int = 'h54f;
    'h186d: romdata_int = 'h1740;
    'h186e: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h186f: romdata_int = 'h55;
    'h1870: romdata_int = 'h6ab;
    'h1871: romdata_int = 'h1156;
    'h1872: romdata_int = 'h421e; // Line descriptor for 1_3s
    'h1873: romdata_int = 'he83;
    'h1874: romdata_int = 'h264;
    'h1875: romdata_int = 'h44c;
    'h1876: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1877: romdata_int = 'he6;
    'h1878: romdata_int = 'h336;
    'h1879: romdata_int = 'habd;
    'h187a: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h187b: romdata_int = 'h18e5;
    'h187c: romdata_int = 'h8b3;
    'h187d: romdata_int = 'h11e;
    'h187e: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h187f: romdata_int = 'h40e;
    'h1880: romdata_int = 'h16a1;
    'h1881: romdata_int = 'h101e;
    'h1882: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1883: romdata_int = 'h832;
    'h1884: romdata_int = 'h441;
    'h1885: romdata_int = 'hd5;
    'h1886: romdata_int = 'h421e; // Line descriptor for 1_3s
    'h1887: romdata_int = 'h722;
    'h1888: romdata_int = 'h8a;
    'h1889: romdata_int = 'h88f;
    'h188a: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h188b: romdata_int = 'h262;
    'h188c: romdata_int = 'h1d13;
    'h188d: romdata_int = 'h1d51;
    'h188e: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h188f: romdata_int = 'h354;
    'h1890: romdata_int = 'h54d;
    'h1891: romdata_int = 'h14a8;
    'h1892: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1893: romdata_int = 'ha5;
    'h1894: romdata_int = 'h8a2;
    'h1895: romdata_int = 'h290;
    'h1896: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1897: romdata_int = 'h8cb;
    'h1898: romdata_int = 'h6b4;
    'h1899: romdata_int = 'hce3;
    'h189a: romdata_int = 'h421e; // Line descriptor for 1_3s
    'h189b: romdata_int = 'h640;
    'h189c: romdata_int = 'hef2;
    'h189d: romdata_int = 'h872;
    'h189e: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h189f: romdata_int = 'h1278;
    'h18a0: romdata_int = 'h698;
    'h18a1: romdata_int = 'h67;
    'h18a2: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h18a3: romdata_int = 'h470;
    'h18a4: romdata_int = 'hcdc;
    'h18a5: romdata_int = 'h618;
    'h18a6: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h18a7: romdata_int = 'h1497;
    'h18a8: romdata_int = 'h8f6;
    'h18a9: romdata_int = 'h538;
    'h18aa: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h18ab: romdata_int = 'h2b6;
    'h18ac: romdata_int = 'h6fd;
    'h18ad: romdata_int = 'he74;
    'h18ae: romdata_int = 'h421e; // Line descriptor for 1_3s
    'h18af: romdata_int = 'hd;
    'h18b0: romdata_int = 'h475;
    'h18b1: romdata_int = 'h8a4;
    'h18b2: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h18b3: romdata_int = 'h1b4d;
    'h18b4: romdata_int = 'h6eb;
    'h18b5: romdata_int = 'h186b;
    'h18b6: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h18b7: romdata_int = 'h2f2;
    'h18b8: romdata_int = 'h1338;
    'h18b9: romdata_int = 'h1a9e;
    'h18ba: romdata_int = 'h221e; // Line descriptor for 1_3s
    'h18bb: romdata_int = 'h128;
    'h18bc: romdata_int = 'h93e;
    'h18bd: romdata_int = 'h1120;
    'h18be: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18bf: romdata_int = 'h6a4;
    'h18c0: romdata_int = 'h80c;
    'h18c1: romdata_int = 'hb67;
    'h18c2: romdata_int = 'h234a;
    'h18c3: romdata_int = 'h431b; // Line descriptor for 2_5s
    'h18c4: romdata_int = 'h2ba;
    'h18c5: romdata_int = 'h68c;
    'h18c6: romdata_int = 'h10ac;
    'h18c7: romdata_int = 'h1cf9;
    'h18c8: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18c9: romdata_int = 'h144;
    'h18ca: romdata_int = 'ha43;
    'h18cb: romdata_int = 'ha74;
    'h18cc: romdata_int = 'h1ac6;
    'h18cd: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18ce: romdata_int = 'h300;
    'h18cf: romdata_int = 'h445;
    'h18d0: romdata_int = 'h451;
    'h18d1: romdata_int = 'h1cd1;
    'h18d2: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18d3: romdata_int = 'h698;
    'h18d4: romdata_int = 'hc35;
    'h18d5: romdata_int = 'h113b;
    'h18d6: romdata_int = 'h20bd;
    'h18d7: romdata_int = 'h431b; // Line descriptor for 2_5s
    'h18d8: romdata_int = 'h8d9;
    'h18d9: romdata_int = 'h924;
    'h18da: romdata_int = 'hc3d;
    'h18db: romdata_int = 'h18b7;
    'h18dc: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18dd: romdata_int = 'h6fc;
    'h18de: romdata_int = 'h54c;
    'h18df: romdata_int = 'h8ed;
    'h18e0: romdata_int = 'h1b54;
    'h18e1: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18e2: romdata_int = 'ha95;
    'h18e3: romdata_int = 'h759;
    'h18e4: romdata_int = 'hd1;
    'h18e5: romdata_int = 'h1911;
    'h18e6: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18e7: romdata_int = 'h4e3;
    'h18e8: romdata_int = 'h89d;
    'h18e9: romdata_int = 'h6d9;
    'h18ea: romdata_int = 'h134c;
    'h18eb: romdata_int = 'h431b; // Line descriptor for 2_5s
    'h18ec: romdata_int = 'h14f4;
    'h18ed: romdata_int = 'ha5d;
    'h18ee: romdata_int = 'h1b;
    'h18ef: romdata_int = 'hef2;
    'h18f0: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18f1: romdata_int = 'h20f;
    'h18f2: romdata_int = 'h2233;
    'h18f3: romdata_int = 'habe;
    'h18f4: romdata_int = 'h100;
    'h18f5: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18f6: romdata_int = 'h1ea4;
    'h18f7: romdata_int = 'h23e;
    'h18f8: romdata_int = 'h808;
    'h18f9: romdata_int = 'ha47;
    'h18fa: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18fb: romdata_int = 'h41;
    'h18fc: romdata_int = 'h99;
    'h18fd: romdata_int = 'h547;
    'h18fe: romdata_int = 'h12d6;
    'h18ff: romdata_int = 'h431b; // Line descriptor for 2_5s
    'h1900: romdata_int = 'ha52;
    'h1901: romdata_int = 'h260;
    'h1902: romdata_int = 'h653;
    'h1903: romdata_int = 'h168e;
    'h1904: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h1905: romdata_int = 'h447;
    'h1906: romdata_int = 'ha12;
    'h1907: romdata_int = 'h17;
    'h1908: romdata_int = 'h2262;
    'h1909: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h190a: romdata_int = 'h241;
    'h190b: romdata_int = 'h1757;
    'h190c: romdata_int = 'h41c;
    'h190d: romdata_int = 'hb59;
    'h190e: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h190f: romdata_int = 'h15;
    'h1910: romdata_int = 'hf6;
    'h1911: romdata_int = 'h1941;
    'h1912: romdata_int = 'h520;
    'h1913: romdata_int = 'h431b; // Line descriptor for 2_5s
    'h1914: romdata_int = 'h718;
    'h1915: romdata_int = 'h71f;
    'h1916: romdata_int = 'hd2e;
    'h1917: romdata_int = 'h1442;
    'h1918: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h1919: romdata_int = 'hab2;
    'h191a: romdata_int = 'h1695;
    'h191b: romdata_int = 'he7c;
    'h191c: romdata_int = 'h730;
    'h191d: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h191e: romdata_int = 'h215d;
    'h191f: romdata_int = 'h2cf;
    'h1920: romdata_int = 'h946;
    'h1921: romdata_int = 'he8a;
    'h1922: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h1923: romdata_int = 'h8a1;
    'h1924: romdata_int = 'h21f;
    'h1925: romdata_int = 'h1ea6;
    'h1926: romdata_int = 'h442;
    'h1927: romdata_int = 'h431b; // Line descriptor for 2_5s
    'h1928: romdata_int = 'h31;
    'h1929: romdata_int = 'h14a3;
    'h192a: romdata_int = 'h965;
    'h192b: romdata_int = 'h276;
    'h192c: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h192d: romdata_int = 'h420;
    'h192e: romdata_int = 'h50c;
    'h192f: romdata_int = 'h1a49;
    'h1930: romdata_int = 'h8b0;
    'h1931: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h1932: romdata_int = 'h1f39;
    'h1933: romdata_int = 'h6c7;
    'h1934: romdata_int = 'h493;
    'h1935: romdata_int = 'ha1d;
    'h1936: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h1937: romdata_int = 'hf8;
    'h1938: romdata_int = 'h328;
    'h1939: romdata_int = 'h820;
    'h193a: romdata_int = 'h1d4d;
    'h193b: romdata_int = 'h431b; // Line descriptor for 2_5s
    'h193c: romdata_int = 'h746;
    'h193d: romdata_int = 'h12a;
    'h193e: romdata_int = 'h1157;
    'h193f: romdata_int = 'h210f;
    'h1940: romdata_int = 'h231b; // Line descriptor for 2_5s
    'h1941: romdata_int = 'h2d2;
    'h1942: romdata_int = 'h303;
    'h1943: romdata_int = 'h94b;
    'h1944: romdata_int = 'h1311;
    'h1945: romdata_int = 'h219; // Line descriptor for 4_9s
    'h1946: romdata_int = 'ha00;
    'h1947: romdata_int = 'h129a;
    'h1948: romdata_int = 'h268a;
    'h1949: romdata_int = 'h319; // Line descriptor for 4_9s
    'h194a: romdata_int = 'h2eb;
    'h194b: romdata_int = 'h425;
    'h194c: romdata_int = 'h4e4;
    'h194d: romdata_int = 'hc00;
    'h194e: romdata_int = 'h4419; // Line descriptor for 4_9s
    'h194f: romdata_int = 'h8f8;
    'h1950: romdata_int = 'h670;
    'h1951: romdata_int = 'h68f;
    'h1952: romdata_int = 'h1d3b;
    'h1953: romdata_int = 'he00;
    'h1954: romdata_int = 'h319; // Line descriptor for 4_9s
    'h1955: romdata_int = 'h2fd;
    'h1956: romdata_int = 'h850;
    'h1957: romdata_int = 'h1000;
    'h1958: romdata_int = 'h2279;
    'h1959: romdata_int = 'h119; // Line descriptor for 4_9s
    'h195a: romdata_int = 'hfe;
    'h195b: romdata_int = 'h1200;
    'h195c: romdata_int = 'h219; // Line descriptor for 4_9s
    'h195d: romdata_int = 'h1a7b;
    'h195e: romdata_int = 'h1400;
    'h195f: romdata_int = 'hc72;
    'h1960: romdata_int = 'h119; // Line descriptor for 4_9s
    'h1961: romdata_int = 'h1600;
    'h1962: romdata_int = 'h1ab8;
    'h1963: romdata_int = 'h4219; // Line descriptor for 4_9s
    'h1964: romdata_int = 'h48c;
    'h1965: romdata_int = 'h1800;
    'h1966: romdata_int = 'h242a;
    'h1967: romdata_int = 'h319; // Line descriptor for 4_9s
    'h1968: romdata_int = 'h1cb9;
    'h1969: romdata_int = 'hce;
    'h196a: romdata_int = 'h102e;
    'h196b: romdata_int = 'h1a00;
    'h196c: romdata_int = 'h219; // Line descriptor for 4_9s
    'h196d: romdata_int = 'h1e9b;
    'h196e: romdata_int = 'h1c00;
    'h196f: romdata_int = 'hb15;
    'h1970: romdata_int = 'h219; // Line descriptor for 4_9s
    'h1971: romdata_int = 'h82f;
    'h1972: romdata_int = 'h2165;
    'h1973: romdata_int = 'h1e00;
    'h1974: romdata_int = 'h319; // Line descriptor for 4_9s
    'h1975: romdata_int = 'h5f;
    'h1976: romdata_int = 'ha2;
    'h1977: romdata_int = 'h2728;
    'h1978: romdata_int = 'h2000;
    'h1979: romdata_int = 'h4319; // Line descriptor for 4_9s
    'h197a: romdata_int = 'he08;
    'h197b: romdata_int = 'h2200;
    'h197c: romdata_int = 'h2a;
    'h197d: romdata_int = 'h1c;
    'h197e: romdata_int = 'h319; // Line descriptor for 4_9s
    'h197f: romdata_int = 'h461;
    'h1980: romdata_int = 'h832;
    'h1981: romdata_int = 'h2400;
    'h1982: romdata_int = 'h24ef;
    'h1983: romdata_int = 'h319; // Line descriptor for 4_9s
    'h1984: romdata_int = 'h27b;
    'h1985: romdata_int = 'h1089;
    'h1986: romdata_int = 'h221e;
    'h1987: romdata_int = 'h2600;
    'h1988: romdata_int = 'h219; // Line descriptor for 4_9s
    'h1989: romdata_int = 'h47f;
    'h198a: romdata_int = 'h8cd;
    'h198b: romdata_int = 'h140b;
    'h198c: romdata_int = 'h119; // Line descriptor for 4_9s
    'h198d: romdata_int = 'h62b;
    'h198e: romdata_int = 'hc02;
    'h198f: romdata_int = 'h4319; // Line descriptor for 4_9s
    'h1990: romdata_int = 'h8bd;
    'h1991: romdata_int = 'h163a;
    'h1992: romdata_int = 'h1859;
    'h1993: romdata_int = 'h6ba;
    'h1994: romdata_int = 'h219; // Line descriptor for 4_9s
    'h1995: romdata_int = 'h265;
    'h1996: romdata_int = 'h493;
    'h1997: romdata_int = 'h1f12;
    'h1998: romdata_int = 'h119; // Line descriptor for 4_9s
    'h1999: romdata_int = 'hf0b;
    'h199a: romdata_int = 'h40a;
    'h199b: romdata_int = 'h319; // Line descriptor for 4_9s
    'h199c: romdata_int = 'h0;
    'h199d: romdata_int = 'hc9;
    'h199e: romdata_int = 'h6b4;
    'h199f: romdata_int = 'h1938;
    'h19a0: romdata_int = 'h219; // Line descriptor for 4_9s
    'h19a1: romdata_int = 'h200;
    'h19a2: romdata_int = 'haa1;
    'h19a3: romdata_int = 'h20c7;
    'h19a4: romdata_int = 'h4319; // Line descriptor for 4_9s
    'h19a5: romdata_int = 'h903;
    'h19a6: romdata_int = 'h400;
    'h19a7: romdata_int = 'h2c0;
    'h19a8: romdata_int = 'h12b0;
    'h19a9: romdata_int = 'h219; // Line descriptor for 4_9s
    'h19aa: romdata_int = 'h2e5;
    'h19ab: romdata_int = 'h600;
    'h19ac: romdata_int = 'h25d;
    'h19ad: romdata_int = 'h2419; // Line descriptor for 4_9s
    'h19ae: romdata_int = 'h16a1;
    'h19af: romdata_int = 'h14ec;
    'h19b0: romdata_int = 'h800;
    'h19b1: romdata_int = 'h6b1;
    'h19b2: romdata_int = 'h6d4;
    'h19b3: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h19b4: romdata_int = 'h165;
    'h19b5: romdata_int = 'h4ac;
    'h19b6: romdata_int = 'h6ee;
    'h19b7: romdata_int = 'hcd4;
    'h19b8: romdata_int = 'h1016;
    'h19b9: romdata_int = 'h1077;
    'h19ba: romdata_int = 'h1200;
    'h19bb: romdata_int = 'h168b;
    'h19bc: romdata_int = 'h250f;
    'h19bd: romdata_int = 'h812; // Line descriptor for 3_5s
    'h19be: romdata_int = 'h313;
    'h19bf: romdata_int = 'h567;
    'h19c0: romdata_int = 'h854;
    'h19c1: romdata_int = 'ha6f;
    'h19c2: romdata_int = 'hd42;
    'h19c3: romdata_int = 'h10e2;
    'h19c4: romdata_int = 'h1278;
    'h19c5: romdata_int = 'h1400;
    'h19c6: romdata_int = 'h34e8;
    'h19c7: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h19c8: romdata_int = 'h216;
    'h19c9: romdata_int = 'h4df;
    'h19ca: romdata_int = 'h55f;
    'h19cb: romdata_int = 'hc5a;
    'h19cc: romdata_int = 'h1031;
    'h19cd: romdata_int = 'h113a;
    'h19ce: romdata_int = 'h1600;
    'h19cf: romdata_int = 'h2035;
    'h19d0: romdata_int = 'h32fd;
    'h19d1: romdata_int = 'h812; // Line descriptor for 3_5s
    'h19d2: romdata_int = 'h228;
    'h19d3: romdata_int = 'h337;
    'h19d4: romdata_int = 'h43e;
    'h19d5: romdata_int = 'h958;
    'h19d6: romdata_int = 'haab;
    'h19d7: romdata_int = 'hb47;
    'h19d8: romdata_int = 'h1451;
    'h19d9: romdata_int = 'h1800;
    'h19da: romdata_int = 'h2cea;
    'h19db: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h19dc: romdata_int = 'h1e;
    'h19dd: romdata_int = 'h79;
    'h19de: romdata_int = 'h245;
    'h19df: romdata_int = 'h109d;
    'h19e0: romdata_int = 'h1063;
    'h19e1: romdata_int = 'h1107;
    'h19e2: romdata_int = 'h1a00;
    'h19e3: romdata_int = 'h233c;
    'h19e4: romdata_int = 'h30bc;
    'h19e5: romdata_int = 'h812; // Line descriptor for 3_5s
    'h19e6: romdata_int = 'h10b;
    'h19e7: romdata_int = 'h291;
    'h19e8: romdata_int = 'h61f;
    'h19e9: romdata_int = 'h708;
    'h19ea: romdata_int = 'h803;
    'h19eb: romdata_int = 'he3e;
    'h19ec: romdata_int = 'h1c00;
    'h19ed: romdata_int = 'h1c60;
    'h19ee: romdata_int = 'h2aa1;
    'h19ef: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h19f0: romdata_int = 'h4c;
    'h19f1: romdata_int = 'h526;
    'h19f2: romdata_int = 'ha94;
    'h19f3: romdata_int = 'haf2;
    'h19f4: romdata_int = 'he79;
    'h19f5: romdata_int = 'h104b;
    'h19f6: romdata_int = 'h1e00;
    'h19f7: romdata_int = 'h1ed2;
    'h19f8: romdata_int = 'h2f21;
    'h19f9: romdata_int = 'h812; // Line descriptor for 3_5s
    'h19fa: romdata_int = 'h13d;
    'h19fb: romdata_int = 'h512;
    'h19fc: romdata_int = 'h6af;
    'h19fd: romdata_int = 'h8e9;
    'h19fe: romdata_int = 'hc2d;
    'h19ff: romdata_int = 'hc80;
    'h1a00: romdata_int = 'h1293;
    'h1a01: romdata_int = 'h2000;
    'h1a02: romdata_int = 'h26b4;
    'h1a03: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h1a04: romdata_int = 'hef;
    'h1a05: romdata_int = 'had3;
    'h1a06: romdata_int = 'hca1;
    'h1a07: romdata_int = 'hd32;
    'h1a08: romdata_int = 'hf0f;
    'h1a09: romdata_int = 'hf39;
    'h1a0a: romdata_int = 'h20ee;
    'h1a0b: romdata_int = 'h2200;
    'h1a0c: romdata_int = 'h2ac7;
    'h1a0d: romdata_int = 'h812; // Line descriptor for 3_5s
    'h1a0e: romdata_int = 'h6e7;
    'h1a0f: romdata_int = 'h8a6;
    'h1a10: romdata_int = 'h8d3;
    'h1a11: romdata_int = 'hb1d;
    'h1a12: romdata_int = 'hb2c;
    'h1a13: romdata_int = 'hcb6;
    'h1a14: romdata_int = 'h1b4c;
    'h1a15: romdata_int = 'h2400;
    'h1a16: romdata_int = 'h2f05;
    'h1a17: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h1a18: romdata_int = 'hbc;
    'h1a19: romdata_int = 'h55a;
    'h1a1a: romdata_int = 'h6bd;
    'h1a1b: romdata_int = 'h8f8;
    'h1a1c: romdata_int = 'hacf;
    'h1a1d: romdata_int = 'hf4e;
    'h1a1e: romdata_int = 'h1e6b;
    'h1a1f: romdata_int = 'h2600;
    'h1a20: romdata_int = 'h2c8e;
    'h1a21: romdata_int = 'h812; // Line descriptor for 3_5s
    'h1a22: romdata_int = 'h99;
    'h1a23: romdata_int = 'h672;
    'h1a24: romdata_int = 'h687;
    'h1a25: romdata_int = 'h85f;
    'h1a26: romdata_int = 'hc30;
    'h1a27: romdata_int = 'he81;
    'h1a28: romdata_int = 'h18dc;
    'h1a29: romdata_int = 'h2800;
    'h1a2a: romdata_int = 'h2908;
    'h1a2b: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h1a2c: romdata_int = 'h27a;
    'h1a2d: romdata_int = 'h2a2;
    'h1a2e: romdata_int = 'h40b;
    'h1a2f: romdata_int = 'h73a;
    'h1a30: romdata_int = 'hb62;
    'h1a31: romdata_int = 'he66;
    'h1a32: romdata_int = 'h144c;
    'h1a33: romdata_int = 'h2a00;
    'h1a34: romdata_int = 'h3510;
    'h1a35: romdata_int = 'h812; // Line descriptor for 3_5s
    'h1a36: romdata_int = 'h20b;
    'h1a37: romdata_int = 'h20e;
    'h1a38: romdata_int = 'hb42;
    'h1a39: romdata_int = 'he5e;
    'h1a3a: romdata_int = 'hec7;
    'h1a3b: romdata_int = 'h10d9;
    'h1a3c: romdata_int = 'h183a;
    'h1a3d: romdata_int = 'h28da;
    'h1a3e: romdata_int = 'h2c00;
    'h1a3f: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h1a40: romdata_int = 'h9d;
    'h1a41: romdata_int = 'hc7;
    'h1a42: romdata_int = 'h506;
    'h1a43: romdata_int = 'h6db;
    'h1a44: romdata_int = 'h817;
    'h1a45: romdata_int = 'heeb;
    'h1a46: romdata_int = 'h1b50;
    'h1a47: romdata_int = 'h240e;
    'h1a48: romdata_int = 'h2e00;
    'h1a49: romdata_int = 'h812; // Line descriptor for 3_5s
    'h1a4a: romdata_int = 'h2a;
    'h1a4b: romdata_int = 'h33e;
    'h1a4c: romdata_int = 'h74f;
    'h1a4d: romdata_int = 'hc45;
    'h1a4e: romdata_int = 'hcc4;
    'h1a4f: romdata_int = 'hf2c;
    'h1a50: romdata_int = 'h22bd;
    'h1a51: romdata_int = 'h3000;
    'h1a52: romdata_int = 'h331b;
    'h1a53: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h1a54: romdata_int = 'h4ed;
    'h1a55: romdata_int = 'h75f;
    'h1a56: romdata_int = 'h886;
    'h1a57: romdata_int = 'h828;
    'h1a58: romdata_int = 'h906;
    'h1a59: romdata_int = 'hafb;
    'h1a5a: romdata_int = 'h1d4e;
    'h1a5b: romdata_int = 'h30da;
    'h1a5c: romdata_int = 'h3200;
    'h1a5d: romdata_int = 'h2812; // Line descriptor for 3_5s
    'h1a5e: romdata_int = 'h34c;
    'h1a5f: romdata_int = 'h540;
    'h1a60: romdata_int = 'hc42;
    'h1a61: romdata_int = 'he0f;
    'h1a62: romdata_int = 'h1047;
    'h1a63: romdata_int = 'h10a3;
    'h1a64: romdata_int = 'h16cd;
    'h1a65: romdata_int = 'h2710;
    'h1a66: romdata_int = 'h3400;
    'h1a67: romdata_int = 'h470f; // Line descriptor for 2_3s
    'h1a68: romdata_int = 'h0;
    'h1a69: romdata_int = 'h134;
    'h1a6a: romdata_int = 'h2c0;
    'h1a6b: romdata_int = 'h162f;
    'h1a6c: romdata_int = 'h16bd;
    'h1a6d: romdata_int = 'h1e00;
    'h1a6e: romdata_int = 'h2443;
    'h1a6f: romdata_int = 'h2e68;
    'h1a70: romdata_int = 'h70f; // Line descriptor for 2_3s
    'h1a71: romdata_int = 'hd5;
    'h1a72: romdata_int = 'he6;
    'h1a73: romdata_int = 'h200;
    'h1a74: romdata_int = 'h265;
    'h1a75: romdata_int = 'h1533;
    'h1a76: romdata_int = 'h1ea9;
    'h1a77: romdata_int = 'h2000;
    'h1a78: romdata_int = 'h2c0f;
    'h1a79: romdata_int = 'h470f; // Line descriptor for 2_3s
    'h1a7a: romdata_int = 'h208;
    'h1a7b: romdata_int = 'h27b;
    'h1a7c: romdata_int = 'h400;
    'h1a7d: romdata_int = 'h407;
    'h1a7e: romdata_int = 'h88f;
    'h1a7f: romdata_int = 'h2200;
    'h1a80: romdata_int = 'h2755;
    'h1a81: romdata_int = 'h2a17;
    'h1a82: romdata_int = 'h70f; // Line descriptor for 2_3s
    'h1a83: romdata_int = 'h67;
    'h1a84: romdata_int = 'h2cf;
    'h1a85: romdata_int = 'h600;
    'h1a86: romdata_int = 'he10;
    'h1a87: romdata_int = 'h1c74;
    'h1a88: romdata_int = 'h20ac;
    'h1a89: romdata_int = 'h2400;
    'h1a8a: romdata_int = 'h32c3;
    'h1a8b: romdata_int = 'h470f; // Line descriptor for 2_3s
    'h1a8c: romdata_int = 'h2eb;
    'h1a8d: romdata_int = 'h2fd;
    'h1a8e: romdata_int = 'h411;
    'h1a8f: romdata_int = 'h6eb;
    'h1a90: romdata_int = 'h800;
    'h1a91: romdata_int = 'h2600;
    'h1a92: romdata_int = 'h3870;
    'h1a93: romdata_int = 'h3a4b;
    'h1a94: romdata_int = 'h70f; // Line descriptor for 2_3s
    'h1a95: romdata_int = 'h61;
    'h1a96: romdata_int = 'h4d0;
    'h1a97: romdata_int = 'ha00;
    'h1a98: romdata_int = 'ha7d;
    'h1a99: romdata_int = 'hd47;
    'h1a9a: romdata_int = 'h2800;
    'h1a9b: romdata_int = 'h306d;
    'h1a9c: romdata_int = 'h362a;
    'h1a9d: romdata_int = 'h470f; // Line descriptor for 2_3s
    'h1a9e: romdata_int = 'ha5;
    'h1a9f: romdata_int = 'h50a;
    'h1aa0: romdata_int = 'hb42;
    'h1aa1: romdata_int = 'hc00;
    'h1aa2: romdata_int = 'h18e4;
    'h1aa3: romdata_int = 'h2a00;
    'h1aa4: romdata_int = 'h2d1e;
    'h1aa5: romdata_int = 'h380f;
    'h1aa6: romdata_int = 'h70f; // Line descriptor for 2_3s
    'h1aa7: romdata_int = 'h11e;
    'h1aa8: romdata_int = 'h560;
    'h1aa9: romdata_int = 'he00;
    'h1aaa: romdata_int = 'h1290;
    'h1aab: romdata_int = 'h12a7;
    'h1aac: romdata_int = 'h275b;
    'h1aad: romdata_int = 'h2c00;
    'h1aae: romdata_int = 'h2e20;
    'h1aaf: romdata_int = 'h470f; // Line descriptor for 2_3s
    'h1ab0: romdata_int = 'h6b;
    'h1ab1: romdata_int = 'h322;
    'h1ab2: romdata_int = 'h4ff;
    'h1ab3: romdata_int = 'h1000;
    'h1ab4: romdata_int = 'h1b00;
    'h1ab5: romdata_int = 'h2526;
    'h1ab6: romdata_int = 'h2e00;
    'h1ab7: romdata_int = 'h3425;
    'h1ab8: romdata_int = 'h70f; // Line descriptor for 2_3s
    'h1ab9: romdata_int = 'he0;
    'h1aba: romdata_int = 'h439;
    'h1abb: romdata_int = 'h4e2;
    'h1abc: romdata_int = 'hd01;
    'h1abd: romdata_int = 'h1200;
    'h1abe: romdata_int = 'h3000;
    'h1abf: romdata_int = 'h349d;
    'h1ac0: romdata_int = 'h3b03;
    'h1ac1: romdata_int = 'h470f; // Line descriptor for 2_3s
    'h1ac2: romdata_int = 'h49c;
    'h1ac3: romdata_int = 'h4b0;
    'h1ac4: romdata_int = 'h1400;
    'h1ac5: romdata_int = 'h189d;
    'h1ac6: romdata_int = 'h1c5a;
    'h1ac7: romdata_int = 'h204e;
    'h1ac8: romdata_int = 'h288f;
    'h1ac9: romdata_int = 'h3200;
    'h1aca: romdata_int = 'h70f; // Line descriptor for 2_3s
    'h1acb: romdata_int = 'h55;
    'h1acc: romdata_int = 'h240;
    'h1acd: romdata_int = 'h105f;
    'h1ace: romdata_int = 'h10c8;
    'h1acf: romdata_int = 'h1600;
    'h1ad0: romdata_int = 'h2ab3;
    'h1ad1: romdata_int = 'h3105;
    'h1ad2: romdata_int = 'h3400;
    'h1ad3: romdata_int = 'h470f; // Line descriptor for 2_3s
    'h1ad4: romdata_int = 'hae;
    'h1ad5: romdata_int = 'h25d;
    'h1ad6: romdata_int = 'h616;
    'h1ad7: romdata_int = 'he66;
    'h1ad8: romdata_int = 'h1800;
    'h1ad9: romdata_int = 'h2266;
    'h1ada: romdata_int = 'h28c2;
    'h1adb: romdata_int = 'h3600;
    'h1adc: romdata_int = 'h70f; // Line descriptor for 2_3s
    'h1add: romdata_int = 'h218;
    'h1ade: romdata_int = 'h2e5;
    'h1adf: romdata_int = 'h917;
    'h1ae0: romdata_int = 'h1442;
    'h1ae1: romdata_int = 'h1a00;
    'h1ae2: romdata_int = 'h1e0a;
    'h1ae3: romdata_int = 'h362d;
    'h1ae4: romdata_int = 'h3800;
    'h1ae5: romdata_int = 'h670f; // Line descriptor for 2_3s
    'h1ae6: romdata_int = 'h8a;
    'h1ae7: romdata_int = 'h40a;
    'h1ae8: romdata_int = 'h43d;
    'h1ae9: romdata_int = 'h1aa4;
    'h1aea: romdata_int = 'h1c00;
    'h1aeb: romdata_int = 'h2221;
    'h1aec: romdata_int = 'h3209;
    'h1aed: romdata_int = 'h3a00;
    'h1aee: romdata_int = 'h70c; // Line descriptor for 11_15s
    'h1aef: romdata_int = 'hda;
    'h1af0: romdata_int = 'h1052;
    'h1af1: romdata_int = 'h1200;
    'h1af2: romdata_int = 'h168f;
    'h1af3: romdata_int = 'h180b;
    'h1af4: romdata_int = 'h2a00;
    'h1af5: romdata_int = 'h36d3;
    'h1af6: romdata_int = 'h40ea;
    'h1af7: romdata_int = 'h490c; // Line descriptor for 11_15s
    'h1af8: romdata_int = 'h54;
    'h1af9: romdata_int = 'h96;
    'h1afa: romdata_int = 'h719;
    'h1afb: romdata_int = 'hb58;
    'h1afc: romdata_int = 'h1400;
    'h1afd: romdata_int = 'h22a2;
    'h1afe: romdata_int = 'h2959;
    'h1aff: romdata_int = 'h2c00;
    'h1b00: romdata_int = 'h3053;
    'h1b01: romdata_int = 'h3318;
    'h1b02: romdata_int = 'h80c; // Line descriptor for 11_15s
    'h1b03: romdata_int = 'h2e;
    'h1b04: romdata_int = 'h93f;
    'h1b05: romdata_int = 'he59;
    'h1b06: romdata_int = 'h1600;
    'h1b07: romdata_int = 'h1a35;
    'h1b08: romdata_int = 'h202d;
    'h1b09: romdata_int = 'h2e00;
    'h1b0a: romdata_int = 'h3452;
    'h1b0b: romdata_int = 'h3a6c;
    'h1b0c: romdata_int = 'h460c; // Line descriptor for 11_15s
    'h1b0d: romdata_int = 'h0;
    'h1b0e: romdata_int = 'h14fa;
    'h1b0f: romdata_int = 'h1800;
    'h1b10: romdata_int = 'h1d1f;
    'h1b11: romdata_int = 'h3000;
    'h1b12: romdata_int = 'h3145;
    'h1b13: romdata_int = 'h3c33;
    'h1b14: romdata_int = 'h70c; // Line descriptor for 11_15s
    'h1b15: romdata_int = 'ha0;
    'h1b16: romdata_int = 'h200;
    'h1b17: romdata_int = 'h1a00;
    'h1b18: romdata_int = 'h2422;
    'h1b19: romdata_int = 'h24a2;
    'h1b1a: romdata_int = 'h3200;
    'h1b1b: romdata_int = 'h3e89;
    'h1b1c: romdata_int = 'h3f03;
    'h1b1d: romdata_int = 'h4a0c; // Line descriptor for 11_15s
    'h1b1e: romdata_int = 'h7b;
    'h1b1f: romdata_int = 'h11e;
    'h1b20: romdata_int = 'h2df;
    'h1b21: romdata_int = 'h400;
    'h1b22: romdata_int = 'h91f;
    'h1b23: romdata_int = 'h1936;
    'h1b24: romdata_int = 'h1a97;
    'h1b25: romdata_int = 'h1c00;
    'h1b26: romdata_int = 'h2e3b;
    'h1b27: romdata_int = 'h3400;
    'h1b28: romdata_int = 'h38c8;
    'h1b29: romdata_int = 'h80c; // Line descriptor for 11_15s
    'h1b2a: romdata_int = 'h10a;
    'h1b2b: romdata_int = 'h600;
    'h1b2c: romdata_int = 'hce4;
    'h1b2d: romdata_int = 'h1279;
    'h1b2e: romdata_int = 'h1e00;
    'h1b2f: romdata_int = 'h26ba;
    'h1b30: romdata_int = 'h345c;
    'h1b31: romdata_int = 'h3600;
    'h1b32: romdata_int = 'h3c0e;
    'h1b33: romdata_int = 'h490c; // Line descriptor for 11_15s
    'h1b34: romdata_int = 'h15e;
    'h1b35: romdata_int = 'h54f;
    'h1b36: romdata_int = 'h800;
    'h1b37: romdata_int = 'h10ba;
    'h1b38: romdata_int = 'h12fc;
    'h1b39: romdata_int = 'h2000;
    'h1b3a: romdata_int = 'h2254;
    'h1b3b: romdata_int = 'h2b00;
    'h1b3c: romdata_int = 'h32c1;
    'h1b3d: romdata_int = 'h3800;
    'h1b3e: romdata_int = 'h80c; // Line descriptor for 11_15s
    'h1b3f: romdata_int = 'ha00;
    'h1b40: romdata_int = 'haab;
    'h1b41: romdata_int = 'hd5c;
    'h1b42: romdata_int = 'h146e;
    'h1b43: romdata_int = 'h1f2e;
    'h1b44: romdata_int = 'h2200;
    'h1b45: romdata_int = 'h2ace;
    'h1b46: romdata_int = 'h2c5a;
    'h1b47: romdata_int = 'h3a00;
    'h1b48: romdata_int = 'h470c; // Line descriptor for 11_15s
    'h1b49: romdata_int = 'h6db;
    'h1b4a: romdata_int = 'hc00;
    'h1b4b: romdata_int = 'h165e;
    'h1b4c: romdata_int = 'h1e68;
    'h1b4d: romdata_int = 'h2400;
    'h1b4e: romdata_int = 'h2cfb;
    'h1b4f: romdata_int = 'h3a9c;
    'h1b50: romdata_int = 'h3c00;
    'h1b51: romdata_int = 'h80c; // Line descriptor for 11_15s
    'h1b52: romdata_int = 'h27;
    'h1b53: romdata_int = 'he00;
    'h1b54: romdata_int = 'hf48;
    'h1b55: romdata_int = 'h1c93;
    'h1b56: romdata_int = 'h2133;
    'h1b57: romdata_int = 'h2600;
    'h1b58: romdata_int = 'h360b;
    'h1b59: romdata_int = 'h388c;
    'h1b5a: romdata_int = 'h3e00;
    'h1b5b: romdata_int = 'h690c; // Line descriptor for 11_15s
    'h1b5c: romdata_int = 'h38;
    'h1b5d: romdata_int = 'h2b1;
    'h1b5e: romdata_int = 'h502;
    'h1b5f: romdata_int = 'h1000;
    'h1b60: romdata_int = 'h2652;
    'h1b61: romdata_int = 'h2800;
    'h1b62: romdata_int = 'h289e;
    'h1b63: romdata_int = 'h2e72;
    'h1b64: romdata_int = 'h4000;
    'h1b65: romdata_int = 'h4075;
    'h1b66: romdata_int = 'h90a; // Line descriptor for 7_9s
    'h1b67: romdata_int = 'h541;
    'h1b68: romdata_int = 'ha00;
    'h1b69: romdata_int = 'hc17;
    'h1b6a: romdata_int = 'h14d3;
    'h1b6b: romdata_int = 'h1e00;
    'h1b6c: romdata_int = 'h20b4;
    'h1b6d: romdata_int = 'h2148;
    'h1b6e: romdata_int = 'h3200;
    'h1b6f: romdata_int = 'h36a1;
    'h1b70: romdata_int = 'h3f5a;
    'h1b71: romdata_int = 'h480a; // Line descriptor for 7_9s
    'h1b72: romdata_int = 'hc00;
    'h1b73: romdata_int = 'h185f;
    'h1b74: romdata_int = 'h1c8e;
    'h1b75: romdata_int = 'h2000;
    'h1b76: romdata_int = 'h2221;
    'h1b77: romdata_int = 'h2c0c;
    'h1b78: romdata_int = 'h3400;
    'h1b79: romdata_int = 'h34bc;
    'h1b7a: romdata_int = 'h370e;
    'h1b7b: romdata_int = 'ha0a; // Line descriptor for 7_9s
    'h1b7c: romdata_int = 'h415;
    'h1b7d: romdata_int = 'h83d;
    'h1b7e: romdata_int = 'he00;
    'h1b7f: romdata_int = 'h1256;
    'h1b80: romdata_int = 'h1b62;
    'h1b81: romdata_int = 'h1ee3;
    'h1b82: romdata_int = 'h2200;
    'h1b83: romdata_int = 'h24ff;
    'h1b84: romdata_int = 'h3248;
    'h1b85: romdata_int = 'h3600;
    'h1b86: romdata_int = 'h38ad;
    'h1b87: romdata_int = 'h490a; // Line descriptor for 7_9s
    'h1b88: romdata_int = 'h2f9;
    'h1b89: romdata_int = 'hb0a;
    'h1b8a: romdata_int = 'h1000;
    'h1b8b: romdata_int = 'h101c;
    'h1b8c: romdata_int = 'h2400;
    'h1b8d: romdata_int = 'h2822;
    'h1b8e: romdata_int = 'h288a;
    'h1b8f: romdata_int = 'h3800;
    'h1b90: romdata_int = 'h3948;
    'h1b91: romdata_int = 'h3c18;
    'h1b92: romdata_int = 'h90a; // Line descriptor for 7_9s
    'h1b93: romdata_int = 'h212;
    'h1b94: romdata_int = 'hf17;
    'h1b95: romdata_int = 'h1200;
    'h1b96: romdata_int = 'h16cb;
    'h1b97: romdata_int = 'h2600;
    'h1b98: romdata_int = 'h2a09;
    'h1b99: romdata_int = 'h2f15;
    'h1b9a: romdata_int = 'h329e;
    'h1b9b: romdata_int = 'h3a00;
    'h1b9c: romdata_int = 'h3d33;
    'h1b9d: romdata_int = 'h4a0a; // Line descriptor for 7_9s
    'h1b9e: romdata_int = 'h0;
    'h1b9f: romdata_int = 'h9c;
    'h1ba0: romdata_int = 'hd0d;
    'h1ba1: romdata_int = 'heca;
    'h1ba2: romdata_int = 'h1400;
    'h1ba3: romdata_int = 'h242e;
    'h1ba4: romdata_int = 'h2800;
    'h1ba5: romdata_int = 'h30b9;
    'h1ba6: romdata_int = 'h3c00;
    'h1ba7: romdata_int = 'h3e5e;
    'h1ba8: romdata_int = 'h4562;
    'h1ba9: romdata_int = 'h4a0a; // Line descriptor for 7_9s
    'h1baa: romdata_int = 'h59;
    'h1bab: romdata_int = 'h200;
    'h1bac: romdata_int = 'h1425;
    'h1bad: romdata_int = 'h1600;
    'h1bae: romdata_int = 'h16e4;
    'h1baf: romdata_int = 'h2a00;
    'h1bb0: romdata_int = 'h2a17;
    'h1bb1: romdata_int = 'h30d3;
    'h1bb2: romdata_int = 'h3e00;
    'h1bb3: romdata_int = 'h40ae;
    'h1bb4: romdata_int = 'h4238;
    'h1bb5: romdata_int = 'h4a0a; // Line descriptor for 7_9s
    'h1bb6: romdata_int = 'h400;
    'h1bb7: romdata_int = 'h648;
    'h1bb8: romdata_int = 'hac2;
    'h1bb9: romdata_int = 'h1800;
    'h1bba: romdata_int = 'h1c1e;
    'h1bbb: romdata_int = 'h1e77;
    'h1bbc: romdata_int = 'h2c00;
    'h1bbd: romdata_int = 'h2e95;
    'h1bbe: romdata_int = 'h3514;
    'h1bbf: romdata_int = 'h4000;
    'h1bc0: romdata_int = 'h428e;
    'h1bc1: romdata_int = 'h4a0a; // Line descriptor for 7_9s
    'h1bc2: romdata_int = 'h600;
    'h1bc3: romdata_int = 'h956;
    'h1bc4: romdata_int = 'h18ce;
    'h1bc5: romdata_int = 'h1a00;
    'h1bc6: romdata_int = 'h1b36;
    'h1bc7: romdata_int = 'h22e6;
    'h1bc8: romdata_int = 'h2667;
    'h1bc9: romdata_int = 'h2e00;
    'h1bca: romdata_int = 'h3a10;
    'h1bcb: romdata_int = 'h4200;
    'h1bcc: romdata_int = 'h4474;
    'h1bcd: romdata_int = 'h6a0a; // Line descriptor for 7_9s
    'h1bce: romdata_int = 'h685;
    'h1bcf: romdata_int = 'h800;
    'h1bd0: romdata_int = 'h112f;
    'h1bd1: romdata_int = 'h1320;
    'h1bd2: romdata_int = 'h1c00;
    'h1bd3: romdata_int = 'h26f7;
    'h1bd4: romdata_int = 'h2d05;
    'h1bd5: romdata_int = 'h3000;
    'h1bd6: romdata_int = 'h3a6d;
    'h1bd7: romdata_int = 'h40cc;
    'h1bd8: romdata_int = 'h4400;
    'h1bd9: romdata_int = 'h4d08; // Line descriptor for 37_45s
    'h1bda: romdata_int = 'h11b;
    'h1bdb: romdata_int = 'h499;
    'h1bdc: romdata_int = 'ha00;
    'h1bdd: romdata_int = 'hb08;
    'h1bde: romdata_int = 'h109e;
    'h1bdf: romdata_int = 'h1a00;
    'h1be0: romdata_int = 'h1e8a;
    'h1be1: romdata_int = 'h1ed4;
    'h1be2: romdata_int = 'h2a00;
    'h1be3: romdata_int = 'h2a20;
    'h1be4: romdata_int = 'h3522;
    'h1be5: romdata_int = 'h3a00;
    'h1be6: romdata_int = 'h452b;
    'h1be7: romdata_int = 'h48d5;
    'h1be8: romdata_int = 'h4d08; // Line descriptor for 37_45s
    'h1be9: romdata_int = 'hb9;
    'h1bea: romdata_int = 'h12d;
    'h1beb: romdata_int = 'hc00;
    'h1bec: romdata_int = 'he44;
    'h1bed: romdata_int = 'h180a;
    'h1bee: romdata_int = 'h1c00;
    'h1bef: romdata_int = 'h1c15;
    'h1bf0: romdata_int = 'h263e;
    'h1bf1: romdata_int = 'h2c00;
    'h1bf2: romdata_int = 'h2e9d;
    'h1bf3: romdata_int = 'h3099;
    'h1bf4: romdata_int = 'h3b28;
    'h1bf5: romdata_int = 'h3c00;
    'h1bf6: romdata_int = 'h3c07;
    'h1bf7: romdata_int = 'h4d08; // Line descriptor for 37_45s
    'h1bf8: romdata_int = 'h669;
    'h1bf9: romdata_int = 'h708;
    'h1bfa: romdata_int = 'he00;
    'h1bfb: romdata_int = 'h131a;
    'h1bfc: romdata_int = 'h160e;
    'h1bfd: romdata_int = 'h1e00;
    'h1bfe: romdata_int = 'h20ef;
    'h1bff: romdata_int = 'h22b5;
    'h1c00: romdata_int = 'h2b36;
    'h1c01: romdata_int = 'h2e00;
    'h1c02: romdata_int = 'h2ecf;
    'h1c03: romdata_int = 'h3e00;
    'h1c04: romdata_int = 'h3e83;
    'h1c05: romdata_int = 'h42d9;
    'h1c06: romdata_int = 'h4d08; // Line descriptor for 37_45s
    'h1c07: romdata_int = 'h0;
    'h1c08: romdata_int = 'h3e;
    'h1c09: romdata_int = 'he66;
    'h1c0a: romdata_int = 'h1000;
    'h1c0b: romdata_int = 'h1918;
    'h1c0c: romdata_int = 'h2000;
    'h1c0d: romdata_int = 'h240b;
    'h1c0e: romdata_int = 'h28c5;
    'h1c0f: romdata_int = 'h3000;
    'h1c10: romdata_int = 'h354e;
    'h1c11: romdata_int = 'h3636;
    'h1c12: romdata_int = 'h3c3c;
    'h1c13: romdata_int = 'h4000;
    'h1c14: romdata_int = 'h4614;
    'h1c15: romdata_int = 'h5008; // Line descriptor for 37_45s
    'h1c16: romdata_int = 'h71;
    'h1c17: romdata_int = 'h59;
    'h1c18: romdata_int = 'h139;
    'h1c19: romdata_int = 'h200;
    'h1c1a: romdata_int = 'h81a;
    'h1c1b: romdata_int = 'hd25;
    'h1c1c: romdata_int = 'h1200;
    'h1c1d: romdata_int = 'h1478;
    'h1c1e: romdata_int = 'h2200;
    'h1c1f: romdata_int = 'h2242;
    'h1c20: romdata_int = 'h2716;
    'h1c21: romdata_int = 'h3200;
    'h1c22: romdata_int = 'h327a;
    'h1c23: romdata_int = 'h381c;
    'h1c24: romdata_int = 'h4200;
    'h1c25: romdata_int = 'h4208;
    'h1c26: romdata_int = 'h494a;
    'h1c27: romdata_int = 'h4f08; // Line descriptor for 37_45s
    'h1c28: romdata_int = 'h29;
    'h1c29: romdata_int = 'h15e;
    'h1c2a: romdata_int = 'h400;
    'h1c2b: romdata_int = 'h847;
    'h1c2c: romdata_int = 'h12d4;
    'h1c2d: romdata_int = 'h1400;
    'h1c2e: romdata_int = 'h172d;
    'h1c2f: romdata_int = 'h1a9b;
    'h1c30: romdata_int = 'h1ac5;
    'h1c31: romdata_int = 'h2400;
    'h1c32: romdata_int = 'h2c8b;
    'h1c33: romdata_int = 'h2c9d;
    'h1c34: romdata_int = 'h3400;
    'h1c35: romdata_int = 'h3aeb;
    'h1c36: romdata_int = 'h4400;
    'h1c37: romdata_int = 'h4650;
    'h1c38: romdata_int = 'h5008; // Line descriptor for 37_45s
    'h1c39: romdata_int = 'h9e;
    'h1c3a: romdata_int = 'hd4;
    'h1c3b: romdata_int = 'h2f0;
    'h1c3c: romdata_int = 'h433;
    'h1c3d: romdata_int = 'h600;
    'h1c3e: romdata_int = 'hd1d;
    'h1c3f: romdata_int = 'h1414;
    'h1c40: romdata_int = 'h1600;
    'h1c41: romdata_int = 'h2479;
    'h1c42: romdata_int = 'h2600;
    'h1c43: romdata_int = 'h2922;
    'h1c44: romdata_int = 'h30b8;
    'h1c45: romdata_int = 'h3600;
    'h1c46: romdata_int = 'h369f;
    'h1c47: romdata_int = 'h3e68;
    'h1c48: romdata_int = 'h40f8;
    'h1c49: romdata_int = 'h4600;
    'h1c4a: romdata_int = 'h6e08; // Line descriptor for 37_45s
    'h1c4b: romdata_int = 'h45;
    'h1c4c: romdata_int = 'h331;
    'h1c4d: romdata_int = 'h800;
    'h1c4e: romdata_int = 'hb29;
    'h1c4f: romdata_int = 'h1011;
    'h1c50: romdata_int = 'h1800;
    'h1c51: romdata_int = 'h1c60;
    'h1c52: romdata_int = 'h2161;
    'h1c53: romdata_int = 'h2800;
    'h1c54: romdata_int = 'h3339;
    'h1c55: romdata_int = 'h3800;
    'h1c56: romdata_int = 'h383e;
    'h1c57: romdata_int = 'h4099;
    'h1c58: romdata_int = 'h4476;
    'h1c59: romdata_int = 'h4800;
    'h1c5a: romdata_int = 'h5805; // Line descriptor for 8_9s
    'h1c5b: romdata_int = 'h0;
    'h1c5c: romdata_int = 'ha1;
    'h1c5d: romdata_int = 'h322;
    'h1c5e: romdata_int = 'h879;
    'h1c5f: romdata_int = 'ha00;
    'h1c60: romdata_int = 'h102a;
    'h1c61: romdata_int = 'h10ef;
    'h1c62: romdata_int = 'h1400;
    'h1c63: romdata_int = 'h1aa7;
    'h1c64: romdata_int = 'h1b2c;
    'h1c65: romdata_int = 'h1e00;
    'h1c66: romdata_int = 'h20e7;
    'h1c67: romdata_int = 'h272b;
    'h1c68: romdata_int = 'h2800;
    'h1c69: romdata_int = 'h284d;
    'h1c6a: romdata_int = 'h2ec0;
    'h1c6b: romdata_int = 'h3200;
    'h1c6c: romdata_int = 'h34cb;
    'h1c6d: romdata_int = 'h38ee;
    'h1c6e: romdata_int = 'h3c00;
    'h1c6f: romdata_int = 'h3c7e;
    'h1c70: romdata_int = 'h44e7;
    'h1c71: romdata_int = 'h4600;
    'h1c72: romdata_int = 'h46c8;
    'h1c73: romdata_int = 'h4d2f;
    'h1c74: romdata_int = 'h5805; // Line descriptor for 8_9s
    'h1c75: romdata_int = 'h200;
    'h1c76: romdata_int = 'h55c;
    'h1c77: romdata_int = 'h6a1;
    'h1c78: romdata_int = 'h739;
    'h1c79: romdata_int = 'hab9;
    'h1c7a: romdata_int = 'hc00;
    'h1c7b: romdata_int = 'he1e;
    'h1c7c: romdata_int = 'h1600;
    'h1c7d: romdata_int = 'h1911;
    'h1c7e: romdata_int = 'h1d2b;
    'h1c7f: romdata_int = 'h1ec9;
    'h1c80: romdata_int = 'h1f54;
    'h1c81: romdata_int = 'h2000;
    'h1c82: romdata_int = 'h2a00;
    'h1c83: romdata_int = 'h2a1e;
    'h1c84: romdata_int = 'h3122;
    'h1c85: romdata_int = 'h3400;
    'h1c86: romdata_int = 'h36fc;
    'h1c87: romdata_int = 'h3af9;
    'h1c88: romdata_int = 'h3e00;
    'h1c89: romdata_int = 'h3e54;
    'h1c8a: romdata_int = 'h446f;
    'h1c8b: romdata_int = 'h467e;
    'h1c8c: romdata_int = 'h4800;
    'h1c8d: romdata_int = 'h4c65;
    'h1c8e: romdata_int = 'h5805; // Line descriptor for 8_9s
    'h1c8f: romdata_int = 'h8e;
    'h1c90: romdata_int = 'h30b;
    'h1c91: romdata_int = 'h400;
    'h1c92: romdata_int = 'h860;
    'h1c93: romdata_int = 'hc9b;
    'h1c94: romdata_int = 'he00;
    'h1c95: romdata_int = 'h128a;
    'h1c96: romdata_int = 'h1455;
    'h1c97: romdata_int = 'h1800;
    'h1c98: romdata_int = 'h1c64;
    'h1c99: romdata_int = 'h2013;
    'h1c9a: romdata_int = 'h2200;
    'h1c9b: romdata_int = 'h2283;
    'h1c9c: romdata_int = 'h2a49;
    'h1c9d: romdata_int = 'h2c00;
    'h1c9e: romdata_int = 'h2c28;
    'h1c9f: romdata_int = 'h3358;
    'h1ca0: romdata_int = 'h3600;
    'h1ca1: romdata_int = 'h3b26;
    'h1ca2: romdata_int = 'h4000;
    'h1ca3: romdata_int = 'h424e;
    'h1ca4: romdata_int = 'h4273;
    'h1ca5: romdata_int = 'h4892;
    'h1ca6: romdata_int = 'h4a00;
    'h1ca7: romdata_int = 'h4eea;
    'h1ca8: romdata_int = 'h5805; // Line descriptor for 8_9s
    'h1ca9: romdata_int = 'h137;
    'h1caa: romdata_int = 'h2ae;
    'h1cab: romdata_int = 'h600;
    'h1cac: romdata_int = 'h8b8;
    'h1cad: romdata_int = 'hb3b;
    'h1cae: romdata_int = 'he79;
    'h1caf: romdata_int = 'h1000;
    'h1cb0: romdata_int = 'h1461;
    'h1cb1: romdata_int = 'h16a5;
    'h1cb2: romdata_int = 'h1a00;
    'h1cb3: romdata_int = 'h2318;
    'h1cb4: romdata_int = 'h2400;
    'h1cb5: romdata_int = 'h2522;
    'h1cb6: romdata_int = 'h2d08;
    'h1cb7: romdata_int = 'h2e00;
    'h1cb8: romdata_int = 'h2e3f;
    'h1cb9: romdata_int = 'h32db;
    'h1cba: romdata_int = 'h351d;
    'h1cbb: romdata_int = 'h3800;
    'h1cbc: romdata_int = 'h3c65;
    'h1cbd: romdata_int = 'h40b3;
    'h1cbe: romdata_int = 'h4200;
    'h1cbf: romdata_int = 'h4911;
    'h1cc0: romdata_int = 'h4b09;
    'h1cc1: romdata_int = 'h4c00;
    'h1cc2: romdata_int = 'h7805; // Line descriptor for 8_9s
    'h1cc3: romdata_int = 'h4e1;
    'h1cc4: romdata_int = 'h4ec;
    'h1cc5: romdata_int = 'h63a;
    'h1cc6: romdata_int = 'h800;
    'h1cc7: romdata_int = 'hd12;
    'h1cc8: romdata_int = 'h1200;
    'h1cc9: romdata_int = 'h1328;
    'h1cca: romdata_int = 'h16e0;
    'h1ccb: romdata_int = 'h18ae;
    'h1ccc: romdata_int = 'h1c00;
    'h1ccd: romdata_int = 'h247c;
    'h1cce: romdata_int = 'h2600;
    'h1ccf: romdata_int = 'h2655;
    'h1cd0: romdata_int = 'h28a1;
    'h1cd1: romdata_int = 'h3000;
    'h1cd2: romdata_int = 'h30cf;
    'h1cd3: romdata_int = 'h3738;
    'h1cd4: romdata_int = 'h386c;
    'h1cd5: romdata_int = 'h3a00;
    'h1cd6: romdata_int = 'h3f54;
    'h1cd7: romdata_int = 'h4038;
    'h1cd8: romdata_int = 'h4400;
    'h1cd9: romdata_int = 'h4a41;
    'h1cda: romdata_int = 'h4e00;
    default: romdata_int = 'h4edc;
  endcase
endmodule

//-------------------------------------------------------------------------
//
// File name    :  ldpc_iocontrol.v
// Title        :
//              :
// Purpose      : Variable node holder/message calculator.  Loads llr
//              : data serially
//
// ----------------------------------------------------------------------
// Revision History :
// ----------------------------------------------------------------------
//   Ver  :| Author   :| Mod. Date   :| Changes Made:
//   v1.0  | JTC      :| 2008/07/02  :|
// ----------------------------------------------------------------------
`timescale 1ns/10ps

module ldpc_iocontrol #(
  parameter FOLDFACTOR     = 4,
  parameter LOG2FOLDFACTOR = 2,
  parameter LASTSHIFTWIDTH = 3,
  parameter NUMINSTANCES   = 180
)(
  input clk,
  input rst,

  // start command, completion indicator
  input      start,
  input[4:0] mode,
  input[5:0] iter_limit,
  output     done,

  // common control outputs
  output iteration,
  output first_iteration,
  output disable_vn,
  output disable_cn,

  // control VN's
  output                     we_vnmsg,
  output[7:0]                addr_vn,
  output[LOG2FOLDFACTOR-1:0] addr_vn_lo,

  // control shuffler
  output                     first_half,
  output[1:0]                shift0,
  output[2:0]                shift1,
  output[LASTSHIFTWIDTH-1:0] shift2,

  // control CN's
  output                     cn_we,
  output                     cn_rd,
  output[7:0]                addr_cn,
  output[LOG2FOLDFACTOR-1:0] addr_cn_lo,

  // ROM
  output[12:0]                  romaddr,
  input[8+5+LASTSHIFTWIDTH-1:0] romdata
);

localparam DONT_SHIFT = 0; // useful for debugging

/*********************************
 * State Machine 1               *
 * Controls the decoding process *
 *********************************/
localparam S_IDLE            = 0;
localparam S_PREPDECODE0     = 1;
localparam S_PREPDECODE1     = 2;
localparam S_FETCHCMD0       = 3;
localparam S_FETCHCMD1       = 4;
localparam S_STOREMSG        = 5;
localparam S_STOREPARITYMSG  = 6;
localparam S_STORESHIFTEDPARITY = 7;
localparam S_FINISHPIPE0     = 8;
localparam S_FINISHPIPE1     = 9;
localparam S_FINISHPIPE2     = 10;
localparam S_FINISHPIPE3     = 11;
localparam S_FINISHPIPE4     = 12;
localparam S_FINISHPIPE5     = 13;
localparam S_FINISHPIPE6     = 14;
localparam S_RESTART         = 15;

localparam TURNAROUND_WAITSTATES = 11;

reg[3:0] state;

reg[7:0] cn_count;
reg[7:0] vn_count;
reg[7:0] ta_count;

reg[12:0] romaddr_int;
reg[12:0] start_addr;
reg[12:0] turnaround_addr;
reg[4:0]  group_depth;
reg       turnaround;
reg       turnaround_next;
reg       last_group;
reg       first_group;
reg       last_group_next;
reg       n64k;
reg[7:0]  q;
reg[4:0]  count;
reg[5:0]  iter_count;
reg       done_int;
reg       first_iteration_int;
reg       iteration_int;

reg first_half_int;

reg[3:0] wait_count;

assign romaddr           = romaddr_int;
assign first_iteration   = first_iteration_int;
assign done              = done_int;
assign first_half        = first_half_int;
assign iteration         = iteration_int;

// synchronous state machine
always @( posedge rst, posedge clk )
  if( rst )
  begin
    state               <= S_IDLE;
    done_int            <= 0;
    iter_count          <= 0;
    romaddr_int         <= 0;
    first_iteration_int <= 0;
    iteration_int       <= 0;
    count               <= 0;
    cn_count            <= 0;
    vn_count            <= 0;
    first_half_int      <= 0;
    romaddr_int         <= 0;
    start_addr          <= 0;
    turnaround_addr     <= 0;
    q                   <= 0;
    turnaround          <= 0;
    turnaround_next     <= 0;
    last_group          <= 0;
    first_group         <= 0;
    n64k                <= 0;
    last_group_next     <= 0;
    group_depth         <= 0;
    wait_count          <= 0;
  end
  else
  begin
    // defaults
    done_int <= 0;

    case( state )
    // wait for start to prepare jump to offset, "mode"
    S_IDLE:
    begin
      if( start )
        state <= S_PREPDECODE0;

      romaddr_int      <= 0;
      romaddr_int[4:0] <= mode;

      iter_count    <= iter_limit;
      iteration_int <= 0;

      first_iteration_int <= 1;
      first_half_int      <= 1;
      cn_count            <= 0;
      vn_count            <= 0;
      ta_count            <= 0;

      first_group <= 1;

      done_int <= 1;
    end

    // "mode" is a pointer to a pointer - jump to mode**
    S_PREPDECODE0:
      state <= S_PREPDECODE1;

    S_PREPDECODE1:
    begin
      state <= S_FETCHCMD0;

      n64k <= romdata[16];

      romaddr_int     <= romdata[12:0];
      start_addr      <= romdata[12:0];
      turnaround_addr <= romdata[12:0];
    end

    // interpret code from ROM
    S_FETCHCMD0:
    begin
      state <= S_FETCHCMD1;

      if( n64k )
        vn_count <= 179;
      else
        vn_count <= 44;
    end

    S_FETCHCMD1:
    begin
      state <= S_STORESHIFTEDPARITY;

      romaddr_int <= romaddr_int + 1;

      turnaround  <= romdata[14];
      last_group  <= romdata[13];
      group_depth <= romdata[12:8];
      q           <= romdata[7:0];
      count       <= 0;
    end

    // write shifted set of parity bits
    S_STORESHIFTEDPARITY:
    begin
      state <= S_STOREMSG;

      romaddr_int <= romaddr_int + 1;
      wait_count  <= TURNAROUND_WAITSTATES;
      first_group <= 0;
    end

    // Write messages
    S_STOREMSG:
    begin
      if( count==group_depth )
        state <= S_STOREPARITYMSG;

      romaddr_int <= romaddr_int + (count!=group_depth);

      count    <= count + 1;
      vn_count <= q + cn_count;
    end

    // write parity bits to CN
    S_STOREPARITYMSG:
    begin
      if( last_group || turnaround )
        state <= S_FINISHPIPE0;
      else
        state <= S_STORESHIFTEDPARITY;

      if( !last_group && !turnaround )
      begin
        cn_count    <= cn_count + 1;
        romaddr_int <= romaddr_int + 1;

        turnaround  <= romdata[14];
        last_group  <= romdata[13];
        group_depth <= romdata[12:8];
        q           <= romdata[7:0];
        count       <= 0;
      end
    end

    // need waitstates between phases to let the pipeline clear out
    S_FINISHPIPE0:
    begin
      if( wait_count==0 )
      begin
        if( last_group && (iter_count==0) && !first_half_int )
        begin
          state    <= S_IDLE;
          done_int <= 1;
        end
        else
          state <= S_RESTART;
      end

      wait_count  <= wait_count - 1;

      if( wait_count==0 )
      begin
        turnaround  <= romdata[14];
        last_group  <= romdata[13];
        group_depth <= romdata[12:8];
        q           <= romdata[7:0];
        count       <= 0;

        cn_count    <= ta_count;
        romaddr_int <= turnaround_addr;

        ta_count        <= cn_count    + 1;
        turnaround_addr <= romaddr_int;

        if( last_group && !first_half_int )
        begin
          cn_count            <= 0;
          iteration_int       <= iteration_int ^ ~first_half_int;
          first_iteration_int <= 0;
          romaddr_int         <= start_addr;
          iter_count          <= iter_count - 1;

          ta_count        <= 0;
          turnaround_addr <= start_addr;
        end
      end
    end

    S_RESTART:
    begin
      state <= S_FETCHCMD1;

      if( cn_count==0 )
      begin
        first_group <= 1;
        if( n64k )
          vn_count <= 179;
        else
          vn_count <= 44;
      end

      first_half_int <= ~first_half_int;
    end

    default: ;
    endcase
  end

  // asynchronous portion of state machine
  reg we;
  reg matchpar;
  reg last_step;

  always @( * )
  begin
    // defaults
    we        <= 0;
    matchpar  <= 0;
    last_step <= 0;

    case( state )
      // Write messages
      S_STOREMSG:
        we <= 1;

      // write parity bits to CN's
      S_STOREPARITYMSG:
      begin
        we       <= 1;
        matchpar <= 1;
      end

      // write parity bits to next CN location
      S_STORESHIFTEDPARITY:
      begin
        we <= 1;

        if( first_group )
          last_step <= 1;
        else
          matchpar  <= 1;
      end

      default: ;
    endcase
  end

/********************************
 * State Machine Helper         *
 * Adds delays to we and to the *
 * addresses for vn and cn      *
 ********************************/
// determine undelayed controls
wire[7:0]                  orig_cn_addr;
wire[7:0]                  orig_vn_addr;
wire[5+LASTSHIFTWIDTH-1:0] orig_shiftval;
wire                       orig_we_vnmsg;
wire                       orig_cn_we;
wire                       orig_cn_rd;
wire                       orig_disable;

assign orig_vn_addr  = ( matchpar || last_step ) ? vn_count
                       : romdata[8+5+LASTSHIFTWIDTH-1:5+LASTSHIFTWIDTH];
assign orig_cn_addr  = cn_count;
assign orig_shiftval = DONT_SHIFT                     ? 0 :
                       matchpar                       ? 0 :
                       (first_half_int && last_step)  ? 1 :
                       (~first_half_int && last_step) ? NUMINSTANCES-1 :
                       first_half_int                 ? romdata[5+LASTSHIFTWIDTH-1:0] :
                                                        NUMINSTANCES - romdata[5+LASTSHIFTWIDTH-1:0];
assign orig_we_vnmsg = we & ~first_half_int;
assign orig_cn_we    = we & first_half_int;
assign orig_cn_rd    = we & ~first_half_int;
assign orig_disable  = last_step;

// add delays to compensate for latencies in external modules
localparam LOCAL_DELAY   = 1;  // Local register delays everything by 1
localparam RAM_LATENCY   = 2;  // RAM registers address in and data out
localparam VN_PIPES      = 3;
localparam SHUFFLE_PIPES = 3;
localparam CN_PIPES      = 2;
localparam MAX_PIPES     = VN_PIPES > CN_PIPES ? VN_PIPES : CN_PIPES;

localparam SHUFFLE_PREPSTAGES = 1; // we'll use 1 pipe locally to calculate shift addresses
localparam DISABLE_PREPSTAGES = 1; // disable needs 1 local pipe to sort out upstream/downstream

localparam LATENCY_VN_DEST  = LOCAL_DELAY + RAM_LATENCY + SHUFFLE_PIPES + CN_PIPES;
localparam LATENCY_CN_DEST  = LOCAL_DELAY + RAM_LATENCY + SHUFFLE_PIPES + VN_PIPES;
localparam LATENCY_CNVN_MAX = LOCAL_DELAY + RAM_LATENCY + SHUFFLE_PIPES + MAX_PIPES;

localparam LATENCY_DISABLE_DL = LATENCY_CN_DEST - DISABLE_PREPSTAGES;
localparam LATENCY_DISABLE_UL = LATENCY_VN_DEST - DISABLE_PREPSTAGES;

localparam LATENCY_SHIFTVALS_DL  = LOCAL_DELAY + RAM_LATENCY + VN_PIPES - SHUFFLE_PREPSTAGES;
localparam LATENCY_SHIFTVALS_UL  = LOCAL_DELAY + RAM_LATENCY + CN_PIPES - SHUFFLE_PREPSTAGES;
localparam LATENCY_SHIFTVALS_MAX = LOCAL_DELAY + RAM_LATENCY + MAX_PIPES - SHUFFLE_PREPSTAGES;

// for code neatness, all shift registers are the same length.  Rely on synthesizer to
// remove unused registers
reg[7:0]                  cn_addr_del[0:LATENCY_CNVN_MAX-1];
reg[7:0]                  vn_addr_del[0:LATENCY_CNVN_MAX-1];
reg[5+LASTSHIFTWIDTH-1:0] shiftval_del[0:LATENCY_CNVN_MAX-1];
reg                       we_vnmsg_del[0:LATENCY_CNVN_MAX-1];
reg                       cn_we_del[0:LATENCY_CNVN_MAX-1];
reg                       cn_rd_del[0:LATENCY_CNVN_MAX-1];
reg                       disable_vn_del[0:LATENCY_CNVN_MAX-1];
reg                       disable_cn_del[0:LATENCY_CNVN_MAX-1];

wire[5+LASTSHIFTWIDTH-1:0] shiftval_int;

integer loopvar;

assign we_vnmsg   = we_vnmsg_del[LATENCY_VN_DEST-1];
assign cn_we      = cn_we_del[LATENCY_CN_DEST-1];
assign cn_rd      = cn_rd_del[LATENCY_CN_DEST-1];
assign addr_vn    = vn_addr_del[LATENCY_VN_DEST-1];
assign addr_cn    = cn_addr_del[LATENCY_CN_DEST-1];
assign disable_vn = disable_vn_del[LATENCY_VN_DEST-1];
assign disable_cn = disable_cn_del[LATENCY_CN_DEST-1];

assign shiftval_int = shiftval_del[LATENCY_SHIFTVALS_MAX-1];

always @( posedge rst, posedge clk )
  if( rst )
    for( loopvar=0; loopvar<LATENCY_CNVN_MAX; loopvar=loopvar+1 )
    begin
      cn_addr_del[loopvar]    <= 0;
      vn_addr_del[loopvar]    <= 0;
      shiftval_del[loopvar]   <= 0;
      we_vnmsg_del[loopvar]   <= 0;
      cn_we_del[loopvar]      <= 0;
      cn_rd_del[loopvar]      <= 0;
      disable_vn_del[loopvar] <= 0;
      disable_cn_del[loopvar] <= 0;
    end
  else
  begin
    cn_addr_del[0]    <= orig_cn_addr;
    vn_addr_del[0]    <= orig_vn_addr;
    shiftval_del[0]   <= orig_shiftval;
    we_vnmsg_del[0]   <= orig_we_vnmsg;
    cn_we_del[0]      <= orig_cn_we;
    cn_rd_del[0]      <= orig_cn_rd;
    disable_vn_del[0] <= orig_disable;
    disable_cn_del[0] <= orig_disable;

    for( loopvar=1; loopvar<LATENCY_CNVN_MAX; loopvar=loopvar+1 )
    begin
      cn_addr_del[loopvar]    <= cn_addr_del[loopvar-1];
      vn_addr_del[loopvar]    <= vn_addr_del[loopvar-1];
      shiftval_del[loopvar]   <= shiftval_del[loopvar-1];
      we_vnmsg_del[loopvar]   <= we_vnmsg_del[loopvar-1];
      cn_we_del[loopvar]      <= cn_we_del[loopvar-1];
      cn_rd_del[loopvar]      <= cn_rd_del[loopvar-1];
      disable_vn_del[loopvar] <= disable_vn_del[loopvar-1];
      disable_cn_del[loopvar] <= disable_cn_del[loopvar-1];
    end

    // need some muxes in the middle of the shift registers because of different
    // latencies for upstream and downstream messages
    if( first_half )
    begin
      vn_addr_del[LATENCY_VN_DEST-1]    <= orig_vn_addr;
      we_vnmsg_del[LATENCY_VN_DEST-1]   <= orig_we_vnmsg;
      disable_vn_del[LATENCY_VN_DEST-1] <= orig_disable;
    end
    if( !first_half )
    begin
      cn_addr_del[LATENCY_CN_DEST-1]    <= orig_cn_addr;
      cn_we_del[LATENCY_CN_DEST-1]      <= orig_cn_we;
      cn_rd_del[LATENCY_CN_DEST-1]      <= orig_cn_rd;
      disable_cn_del[LATENCY_CN_DEST-1] <= orig_disable;
    end
    
    if( first_half )
      shiftval_del[LATENCY_SHIFTVALS_MAX-1] <= shiftval_del[LATENCY_SHIFTVALS_DL-2];
    if( !first_half )
      shiftval_del[LATENCY_SHIFTVALS_MAX-1] <= shiftval_del[LATENCY_SHIFTVALS_UL-2];
  end

wire[1:0]               shift0_int;
reg[1:0]                shift0_reg;
wire[2:0]               shift1_int;
reg[2:0]                shift1_reg;
reg[LASTSHIFTWIDTH-1:0] shift2_reg;

assign shift0 = shift0_reg;
assign shift1 = shift1_reg;
assign shift2 = shift2_reg;

reg[8:0]                rem0;
reg[LASTSHIFTWIDTH-1:0] rem1;

generate
  if( FOLDFACTOR==1 )
  begin: case360
    assign shift0_int = shiftval_int > 269 ? 3
                      : shiftval_int > 179 ? 2
                      : shiftval_int > 89  ? 1
                      :                      0;

    assign shift1_int = rem0 > 83 ? 7
                      : rem0 > 71 ? 6
                      : rem0 > 59 ? 5
                      : rem0 > 47 ? 4
                      : rem0 > 35 ? 3
                      : rem0 > 23 ? 2
                      : rem0 > 11 ? 1
                      :             0;
  end
  if( FOLDFACTOR==2 )
  begin: case180
    assign shift0_int = shiftval_int > 134 ? 3
                      : shiftval_int > 89  ? 2
                      : shiftval_int > 44  ? 1
                      :                      0;


    assign shift1_int = rem0 > 41 ? 7
                      : rem0 > 35 ? 6
                      : rem0 > 29 ? 5
                      : rem0 > 23 ? 4
                      : rem0 > 17 ? 3
                      : rem0 > 11 ? 2
                      : rem0 > 5  ? 1
                      :             0;
  end
  if( FOLDFACTOR==3 )
  begin: case120
    assign shift0_int = shiftval_int > 89 ? 3
                      : shiftval_int > 59 ? 2
                      : shiftval_int > 29 ? 1
                      :                     0;

    assign shift1_int = rem0 > 26 ? 7
                      : rem0 > 22 ? 6
                      : rem0 > 18 ? 5
                      : rem0 > 15 ? 4
                      : rem0 > 11 ? 3
                      : rem0 > 7  ? 2
                      : rem0 > 3  ? 1
                      :             0;
  end
  if( FOLDFACTOR==4 )
  begin: case90
    assign shift0_int = shiftval_int > 66 ? 3
                      : shiftval_int > 44 ? 2
                      : shiftval_int > 22 ? 1
                      :                     0;

    assign shift1_int = rem0 > 20 ? 7
                      : rem0 > 17 ? 6
                      : rem0 > 14 ? 5
                      : rem0 > 11 ? 4
                      : rem0 > 8  ? 3
                      : rem0 > 5  ? 2
                      : rem0 > 2  ? 1
                      :             0;
  end
endgenerate

always @( posedge rst, posedge clk )
  if( rst )
  begin
    shift0_reg            <= 0;
    shift1_reg            <= 0;
    shift2_reg            <= 0;
    rem0                  <= 0;
    rem1                  <= 0;
  end
  else
  begin
    // shift0 needs to be inverted (this arithmetic should be optimized out)
    shift0_reg <= shift0_int;
    shift1_reg <= shift1_int;
    shift2_reg <= rem1;

    // calculate remainders after first two shifts
    if( FOLDFACTOR==1 )
      rem0 <= shift0_int==3 ? shiftval_int-270
            : shift0_int==2 ? shiftval_int-180
            : shift0_int==1 ? shiftval_int-90
            :                 shiftval_int;
    if( FOLDFACTOR==2 )
      rem0 <= shift0_int==3 ? shiftval_int-135
            : shift0_int==2 ? shiftval_int-90
            : shift0_int==1 ? shiftval_int-45
            :                 shiftval_int;
    if( FOLDFACTOR==3 )
      rem0 <= shift0_int==3 ? shiftval_int-90
            : shift0_int==2 ? shiftval_int-60
            : shift0_int==1 ? shiftval_int-30
            :                 shiftval_int;
    if( FOLDFACTOR==4 )
      rem0 <= shift0_int==3 ? shiftval_int-67
            : shift0_int==2 ? shiftval_int-45
            : shift0_int==1 ? shiftval_int-23
            :                 shiftval_int;

    if( FOLDFACTOR==1 )
      rem1 <= shift1_int==7 ? rem0-84
            : shift1_int==6 ? rem0-72
            : shift1_int==5 ? rem0-60
            : shift1_int==4 ? rem0-48
            : shift1_int==3 ? rem0-36
            : shift1_int==2 ? rem0-24
            : shift1_int==1 ? rem0-12
            :                 rem0;
    if( FOLDFACTOR==3 )
      rem1 <= shift1_int==7 ? rem0-52
            : shift1_int==6 ? rem0-45
            : shift1_int==5 ? rem0-37
            : shift1_int==4 ? rem0-30
            : shift1_int==3 ? rem0-22
            : shift1_int==2 ? rem0-15
            : shift1_int==1 ? rem0-7
            :                 rem0;
    if( FOLDFACTOR==4 )
      rem1 <= shift1_int==7 ? rem0-21
            : shift1_int==6 ? rem0-18
            : shift1_int==5 ? rem0-15
            : shift1_int==4 ? rem0-12
            : shift1_int==3 ? rem0-9
            : shift1_int==2 ? rem0-6
            : shift1_int==1 ? rem0-3
            :                 rem0;
  end
endmodule
//-------------------------------------------------------------------------
//
// File name    :  ldpc_muxreg.v
// Title        :
//              :
// Purpose      : Just a multiplexer and a register, but I added a level
//              : of hierarchy because design_vision was choking on the
//              : flat version
//
// ----------------------------------------------------------------------
// Revision History :
// ----------------------------------------------------------------------
//   Ver  :| Author   :| Mod. Date   :| Changes Made:
//   v1.0  | JTC      :| 2008/07/02  :|
// ----------------------------------------------------------------------
`timescale 1ns/10ps

module ldpc_muxreg #(
  parameter LLRWIDTH = 4,
  parameter NUMINPS  = 4,
  parameter MUXSIZE  = 4,
  parameter SELBITS  = 2
)(
  input clk,
  input rst,

  input[SELBITS-1:0]          sel,
  input[NUMINPS*LLRWIDTH-1:0] din,
  output[LLRWIDTH-1:0]        dout
);

// convert to 2-d array
wire[LLRWIDTH-1:0] din_2d[MUXSIZE-1:0];

generate
  genvar muxpos;

  for( muxpos=0; muxpos<MUXSIZE; muxpos=muxpos+1 )
  begin: muxto2d
    assign din_2d[muxpos] = din[muxpos*LLRWIDTH+LLRWIDTH-1 -: LLRWIDTH];
  end
endgenerate

// mux and register
reg[LLRWIDTH-1:0] mux_result;

assign dout = mux_result;

always @( posedge clk, posedge rst )
  if( rst )
    mux_result <= 0;
  else
    mux_result <= din_2d[sel];
endmodule
//-------------------------------------------------------------------------
//
// File name    :  ldpc_ram_behav.v
// Title        :
//              :
// Purpose      : RAM behavioral model
//
// ----------------------------------------------------------------------
// Revision History :
// ----------------------------------------------------------------------
//   Ver  :| Author   :| Mod. Date   :| Changes Made:
//   v1.0  | JTC      :| 2008/07/02  :|
// ----------------------------------------------------------------------
`timescale 1ns/10ps

module ldpc_ram_behav #(
  parameter WIDTH     = 4,
  parameter LOG2DEPTH = 4
)(
  input                clk,
  input                we,
  input[WIDTH-1:0]     din,
  input[LOG2DEPTH-1:0] wraddr,
  input[LOG2DEPTH-1:0] rdaddr,
  output[WIDTH-1:0]    dout
);

reg[WIDTH-1:0]     storage[0:2**LOG2DEPTH -1];
reg[LOG2DEPTH-1:0] addr_del;
reg[WIDTH-1:0]     dout_int;

assign dout = dout_int;

always @( posedge clk )
begin
  if( !we )
    storage[wraddr] <= din;
  
  addr_del <= rdaddr;
  
  dout_int <= storage[addr_del];
end

endmodule
//-------------------------------------------------------------------------
//
// File name    :  ldpc_shuffle.v
// Title        :
//              :
// Purpose      : Barrel-rotate of NUINSTANCES, LLRWIDTH-bit inputs
//
// ----------------------------------------------------------------------
// Revision History :
// ----------------------------------------------------------------------
//   Ver  :| Author   :| Mod. Date   :| Changes Made:
//   v1.0  | JTC      :| 2008/07/02  :|
// ----------------------------------------------------------------------
`timescale 1ns/10ps

module ldpc_shuffle #(
  parameter FOLDFACTOR     = 4,
  parameter NUMINSTANCES   = 360/FOLDFACTOR,
  parameter LOG2INSTANCES  = 10 - FOLDFACTOR,
  parameter LLRWIDTH       = 4,
  parameter LASTSHIFTWIDTH = 3,
  parameter LASTSHIFTDIST  = 6
)(
  input clk,
  input rst,

  // control inputs
  input                     first_half,
  input[1:0]                shift0,
  input[2:0]                shift1,
  input[LASTSHIFTWIDTH-1:0] shift2,

  // message I/O
  input[NUMINSTANCES*LLRWIDTH-1:0]  vn_concat,
  input[NUMINSTANCES*LLRWIDTH-1:0]  cn_concat,
  output[NUMINSTANCES*LLRWIDTH-1:0] sh_concat
);

/*----------------*
 * Shift stage 0  *
 *----------------*/
wire[LLRWIDTH-1:0]     unshifted[NUMINSTANCES-1:0];
wire[LLRWIDTH-1:0]     shifted_0[NUMINSTANCES-1:0];

// convert to 2-d array to make simulation easier to follow, and mux vn/cn msgs
generate
  genvar vecpos;

  for( vecpos=0; vecpos<NUMINSTANCES; vecpos=vecpos+1 )
  begin: to2d
    assign unshifted[vecpos] =
      first_half ? vn_concat[vecpos*LLRWIDTH+LLRWIDTH-1 -: LLRWIDTH]
                 : cn_concat[vecpos*LLRWIDTH+LLRWIDTH-1 -: LLRWIDTH];
  end
endgenerate

// shift distance is shift0* SHIFT0_MULT, where SHIFT0_MULT=
// ceiling(360/FOLDFACTOR/4)
localparam SHIFT0_MULT = (FOLDFACTOR==1) ? 90 :
                         (FOLDFACTOR==2) ? 45 :
                         (FOLDFACTOR==3) ? 30 :
                         /* 4 */           23;

generate
  genvar pos0;

  for( pos0=0; pos0<NUMINSTANCES; pos0=pos0+1 )
  begin: quartershift
    wire[4*LLRWIDTH-1:0] muxinp0;

    assign muxinp0 = { unshifted[(NUMINSTANCES+pos0-3*SHIFT0_MULT) %NUMINSTANCES],
                       unshifted[(NUMINSTANCES+pos0-2*SHIFT0_MULT) %NUMINSTANCES],
                       unshifted[(NUMINSTANCES+pos0-  SHIFT0_MULT) %NUMINSTANCES],
                       unshifted[pos0]  };

    ldpc_muxreg #(
      .LLRWIDTH(LLRWIDTH),
      .NUMINPS (4),
      .MUXSIZE (4),
      .SELBITS (2)
    ) ldpc_muxregi (
      .clk( clk ),
      .rst( rst ),
      .sel( shift0 ),
      .din( muxinp0 ),
      .dout( shifted_0[pos0] )
    );
  end
endgenerate

/*----------------*
 * Shift stage 1  *
 *----------------*/
wire[LLRWIDTH-1:0]     shifted_1[NUMINSTANCES-1:0];

// shift distance is shift1* SHIFT1_MULT, where SHIFT1_MULT=
// ceiling(360/FOLDFACTOR/4/8)
localparam SHIFT1_MULT = (FOLDFACTOR==1) ? 12 :
                         (FOLDFACTOR==2) ? 6  :
                         (FOLDFACTOR==3) ? 4  :
                         /* 4 */           3;

generate
  genvar pos1;

  for( pos1=0; pos1<NUMINSTANCES; pos1=pos1+1 )
  begin: middleshift
    wire[8*LLRWIDTH-1:0] muxinp1;

    assign muxinp1 = { shifted_0[(NUMINSTANCES+pos1-7*SHIFT1_MULT) %NUMINSTANCES],
                       shifted_0[(NUMINSTANCES+pos1-6*SHIFT1_MULT) %NUMINSTANCES],
                       shifted_0[(NUMINSTANCES+pos1-5*SHIFT1_MULT) %NUMINSTANCES],
                       shifted_0[(NUMINSTANCES+pos1-4*SHIFT1_MULT) %NUMINSTANCES],
                       shifted_0[(NUMINSTANCES+pos1-3*SHIFT1_MULT) %NUMINSTANCES],
                       shifted_0[(NUMINSTANCES+pos1-2*SHIFT1_MULT) %NUMINSTANCES],
                       shifted_0[(NUMINSTANCES+pos1-  SHIFT1_MULT) %NUMINSTANCES],
                       shifted_0[pos1]  };

    ldpc_muxreg #(
      .LLRWIDTH(LLRWIDTH),
      .NUMINPS (8),
      .MUXSIZE (8),
      .SELBITS (3)
    ) ldpc_muxregi (
      .clk( clk ),
      .rst( rst ),
      .sel( shift1 ),
      .din( muxinp1 ),
      .dout( shifted_1[pos1] )
    );
  end
endgenerate
  
/*----------------*
 * Shift stage 2  *
 *----------------*/
// This stage is a little more complicated than the others, since there is a
// maximum shift distance
wire[LLRWIDTH-1:0]    shifted_2[NUMINSTANCES-1:0];
reg[NUMINSTANCES-1:0] increment_int;

generate
  genvar pos2;

  for( pos2=0; pos2<NUMINSTANCES; pos2=pos2+1 )
  begin: lastshift
    wire[12*LLRWIDTH-1:0] muxinp2;
    
    assign muxinp2 = { shifted_1[(NUMINSTANCES+pos2-11) %NUMINSTANCES],
                       shifted_1[(NUMINSTANCES+pos2-10) %NUMINSTANCES],
                       shifted_1[(NUMINSTANCES+pos2-9)  %NUMINSTANCES],
                       shifted_1[(NUMINSTANCES+pos2-8)  %NUMINSTANCES],
                       shifted_1[(NUMINSTANCES+pos2-7)  %NUMINSTANCES],
                       shifted_1[(NUMINSTANCES+pos2-6)  %NUMINSTANCES],
                       shifted_1[(NUMINSTANCES+pos2-5)  %NUMINSTANCES],
                       shifted_1[(NUMINSTANCES+pos2-4)  %NUMINSTANCES],
                       shifted_1[(NUMINSTANCES+pos2-3)  %NUMINSTANCES],
                       shifted_1[(NUMINSTANCES+pos2-2)  %NUMINSTANCES],
                       shifted_1[(NUMINSTANCES+pos2-1)  %NUMINSTANCES],
                       shifted_1[pos2]  };

    ldpc_muxreg #(
      .LLRWIDTH(LLRWIDTH),
      .NUMINPS (12),
      .MUXSIZE ((LASTSHIFTDIST+1)),
      .SELBITS (LASTSHIFTWIDTH)
    ) ldpc_muxregi (
      .clk( clk ),
      .rst( rst ),
      .sel( shift2 ),
      .din( muxinp2 ),
      .dout( shifted_2[pos2] )
    );
  end
endgenerate

// assign 2-d array to 1-d output port
generate
  genvar ovecpos;

  for( ovecpos=0; ovecpos<NUMINSTANCES; ovecpos=ovecpos+1 )
  begin: to1d
    assign sh_concat[ovecpos*LLRWIDTH+LLRWIDTH-1 -: LLRWIDTH] =
              shifted_2[ovecpos];
  end
endgenerate

// decode
localparam SECTION_LEN = (FOLDFACTOR==1) ? 90 :
                         (FOLDFACTOR==2) ? 45 :
                         (FOLDFACTOR==3) ? 30 :
                                           23;
function[SECTION_LEN-1:0] Decoder( input[LOG2INSTANCES-3:0] incpointxx );
  integer position;
begin
  Decoder[0] = incpointxx==0;
  
  for( position=1; position<SECTION_LEN; position=position+1 )
    Decoder[position] = (incpointxx==position) || Decoder[position-1];
end
endfunction

endmodule
//-------------------------------------------------------------------------
//
// File name    :  ldp_top.v
// Title        :
//              :
// Purpose      : Top-level of LDPC decoder, structural verilog only
//
// ----------------------------------------------------------------------
// Revision History :
// ----------------------------------------------------------------------
//   Ver  :| Author   :| Mod. Date   :| Changes Made:
//   v1.0  | JTC      :| 2008/07/02  :|
// ----------------------------------------------------------------------
`timescale 1ns/10ps

module ldp_top #(
  parameter FOLDFACTOR     = 4,
  parameter LOG2FOLDFACTOR = 2,
  parameter NUMINSTANCES   = 360,
  parameter LLRWIDTH       = 6
)(
  input clk,
  input rst,

  // LLR I/O
  input                             llr_access,
  input[7+FOLDFACTOR-1:0]           llr_addr,
  input                             llr_din_we,
  input[NUMINSTANCES*LLRWIDTH-1:0]  llr_din,
  output[NUMINSTANCES*LLRWIDTH-1:0] llr_dout,

  // start command, completion indicator
  input      start,
  input[4:0] mode,
  input[5:0] iter_limit,
  output     done
);

////////////////
// PARAMETERS //
////////////////
localparam NUMVNS       = 3;
localparam LASTSHIFTDIST = (FOLDFACTOR==1) ? 11 :
                           (FOLDFACTOR==2) ? 5  :
                           (FOLDFACTOR==3) ? 3  :
                           /* 4 */           2;
localparam LASTSHIFTWIDTH  = (FOLDFACTOR==1) ? 4 :
                             (FOLDFACTOR==2) ? 3 :
                             (FOLDFACTOR==3) ? 2 :
                             /* 4 */           2;

//////////////////////
// INTERNAL SIGNALS //
//////////////////////
wire   zero;
assign zero = 0;

// iocontrol common control outputs
wire iteration;
wire first_iteration;
wire disable_vn;
wire disable_cn;

// iocontrol VN controls
wire                   we_vnmsg;
wire[7+FOLDFACTOR-1:0] addr_vn;

// iocontrol shuffler controls
wire                     first_half;
wire[1:0]                shift0;
wire[2:0]                shift1;
wire[LASTSHIFTWIDTH-1:0] shift2;

// iocontrol CN controls
wire                   cn_we;
wire                   cn_rd;
wire[7+FOLDFACTOR-1:0] addr_cn;

// iocontrol ROM
wire[12:0]                   romaddr;
wire[8+5+LASTSHIFTWIDTH-1:0] romdata;

////////////////////
// Control module //
////////////////////
ldpc_iocontrol #(
  .FOLDFACTOR(FOLDFACTOR),
  .LASTSHIFTWIDTH(LASTSHIFTWIDTH),
  .NUMINSTANCES(NUMINSTANCES)
)
ldpc_iocontroli(
  .clk              (clk),
  .rst              (rst),
  
  .start            (start),
  .mode             (mode),
  .iter_limit       (iter_limit),
  .done             (done),
  
  .iteration        (iteration),
  .first_iteration  (first_iteration),
  .disable_vn       (disable_vn),
  .disable_cn       (disable_cn),
  
  .we_vnmsg         (we_vnmsg),
  .addr_vn          (addr_vn),
  .addr_vn_lo       (),
  
  .first_half       (first_half),
  .shift0           (shift0),
  .shift1           (shift1),
  .shift2           (shift2),

  .cn_we            (cn_we),
  .cn_rd            (cn_rd),
  .addr_cn          (addr_cn),
  .addr_cn_lo       (),

  .romaddr          (romaddr),
  .romdata          (romdata)
);

// asynchronous ROM, attached to control module
ldpc_edgetable ldpc_edgetable_i(
  .clk     ( clk ),
  .rst     ( rst ),
  .romaddr ( romaddr ),
  .romdata ( romdata )
);

////////////////////////
// 2-d/1-d conversion //
////////////////////////
wire[NUMINSTANCES*LLRWIDTH-1:0] cn_concat;
wire[LLRWIDTH-1:0] cn_msg[0:NUMINSTANCES-1];
wire[NUMINSTANCES*LLRWIDTH-1:0] sh_concat;
wire[LLRWIDTH-1:0] sh_msg[0:NUMINSTANCES-1];


generate
  genvar j;

  for( j=0; j<NUMINSTANCES; j=j+1 )
  begin: convert1d2d
    assign cn_concat[LLRWIDTH*j+LLRWIDTH-1 -: LLRWIDTH] = cn_msg[j];
    assign sh_msg[j] = sh_concat[LLRWIDTH*j+LLRWIDTH-1 -: LLRWIDTH];
  end
endgenerate

wire[NUMVNS*LLRWIDTH-1:0]       vn_cluster_msg[0:NUMINSTANCES/NUMVNS-1];
wire[NUMINSTANCES*LLRWIDTH-1:0] vn_concat;
wire[NUMVNS*LLRWIDTH-1:0]       sh_cluster_msg[0:NUMINSTANCES/NUMVNS-1];

wire[NUMVNS*LLRWIDTH-1:0] llr_din_2d[0:NUMINSTANCES/NUMVNS-1];
wire[NUMVNS*LLRWIDTH-1:0] llr_dout_2d[0:NUMINSTANCES/NUMVNS-1];

generate
  genvar m;

  for( m=0; m<NUMINSTANCES/NUMVNS; m=m+1 )
  begin: convert1d2d2
    assign vn_concat[NUMVNS*LLRWIDTH*m+NUMVNS*LLRWIDTH-1 -: NUMVNS*LLRWIDTH] = vn_cluster_msg[m];
    assign sh_cluster_msg[m] = sh_concat[NUMVNS*LLRWIDTH*m+NUMVNS*LLRWIDTH-1 -: NUMVNS*LLRWIDTH];

    assign llr_din_2d[m] = llr_din[NUMVNS*LLRWIDTH*m+NUMVNS*LLRWIDTH-1 -: NUMVNS*LLRWIDTH];
    assign llr_dout[NUMVNS*LLRWIDTH*m+NUMVNS*LLRWIDTH-1 -: NUMVNS*LLRWIDTH] = llr_dout_2d[m];
  end
endgenerate

//////////
// VN's //
//////////
generate
  genvar i;

  for( i=0; i<NUMINSTANCES/NUMVNS; i=i+1 )
  begin: varnodes
    // first
    if( i==0 )
    begin
      ldpc_vncluster #(
        .NUMVNS         (NUMVNS),
        .ENABLE_DISABLE (0),
        .FOLDFACTOR     (FOLDFACTOR),
        .LASTSHIFTWIDTH (LASTSHIFTWIDTH),
        .LLRWIDTH       (LLRWIDTH)
      ) ldpc_vncluster_firsti(
        .clk              (clk),
        .rst              (rst),
        .llr_access       (llr_access),
        .llr_addr         (llr_addr),
        .llr_din_we       (llr_din_we),
        .llr_din          (llr_din_2d[i]),
        .llr_dout         (llr_dout_2d[i]),
        .iteration        (iteration),
        .first_half       (first_half),
        .first_iteration  (first_iteration),
        .we_vnmsg         (we_vnmsg),
        .disable_vn       (zero),
        .addr_vn          (addr_vn),
        .sh_cluster_msg     (sh_cluster_msg[i]),
        .vn_cluster_msg     (vn_cluster_msg[i])
      );
    end

    // last
    if( i==NUMINSTANCES/NUMVNS-1 )
    begin
      ldpc_vncluster #(
        .NUMVNS         (NUMVNS),
        .ENABLE_DISABLE (1),
        .FOLDFACTOR     (FOLDFACTOR),
        .LASTSHIFTWIDTH (LASTSHIFTWIDTH),
        .LLRWIDTH       (LLRWIDTH)
      ) ldpc_vncluster_lasti(
        .clk              (clk),
        .rst              (rst),
        .llr_access       (llr_access),
        .llr_addr         (llr_addr),
        .llr_din_we       (llr_din_we),
        .llr_din          (llr_din_2d[i]),
        .llr_dout         (llr_dout_2d[i]),
        .iteration        (iteration),
        .first_half       (first_half),
        .first_iteration  (first_iteration),
        .we_vnmsg         (we_vnmsg),
        .disable_vn       (disable_vn),
        .addr_vn          (addr_vn),
        .sh_cluster_msg   (sh_cluster_msg[i]),
        .vn_cluster_msg   (vn_cluster_msg[i])
      );
    end

    if( (i!=0) && (i!=NUMINSTANCES/NUMVNS-1) )
    begin
      ldpc_vncluster #(
        .NUMVNS         (NUMVNS),
        .ENABLE_DISABLE (0),
        .FOLDFACTOR     (FOLDFACTOR),
        .LASTSHIFTWIDTH (LASTSHIFTWIDTH),
        .LLRWIDTH       (LLRWIDTH)
      ) ldpc_vnclusteri(
        .clk              (clk),
        .rst              (rst),
        .llr_access       (llr_access),
        .llr_addr         (llr_addr),
        .llr_din_we       (llr_din_we),
        .llr_din          (llr_din_2d[i]),
        .llr_dout         (llr_dout_2d[i]),
        .iteration        (iteration),
        .first_half       (first_half),
        .first_iteration  (first_iteration),
        .we_vnmsg         (we_vnmsg),
        .disable_vn       (zero),
        .addr_vn          (addr_vn),
        .sh_cluster_msg   (sh_cluster_msg[i]),
        .vn_cluster_msg   (vn_cluster_msg[i])
      );
    end
  end
endgenerate

//////////////
// SHUFFLER //
//////////////
ldpc_shuffle #( .FOLDFACTOR(FOLDFACTOR),
                .NUMINSTANCES(NUMINSTANCES),
                .LLRWIDTH(LLRWIDTH),
                .LASTSHIFTWIDTH(LASTSHIFTWIDTH),
                .LASTSHIFTDIST(LASTSHIFTDIST)
 ) ldpc_shufflei(
  .clk          (clk),
  .rst          (rst),
  .first_half   (first_half),
  .shift0       (shift0),
  .shift1       (shift1),
  .shift2       (shift2),
  .vn_concat    (vn_concat),
  .cn_concat    (cn_concat),
  .sh_concat    (sh_concat)
);

//////////
// CN's //
//////////
wire                         dnmsg_we;
wire                         dnmsg_we_gated;
wire[7+FOLDFACTOR-1:0]       dnmsg_wraddr[0:NUMINSTANCES-1];
wire[7+FOLDFACTOR-1:0]       dnmsg_rdaddr[0:NUMINSTANCES-1];
wire[17+4*(LLRWIDTH-1)+31:0] dnmsg_din[0:NUMINSTANCES-1];
wire[17+4*(LLRWIDTH-1)+31:0] dnmsg_dout[0:NUMINSTANCES-1];

// first
ldpc_cn #( .FOLDFACTOR(FOLDFACTOR),
           .LLRWIDTH(LLRWIDTH)
) ldpc_cn0i(
  .clk              (clk),
  .rst              (rst),
  .llr_access       (llr_access),
  .llr_addr         (llr_addr),
  .llr_din_we       (llr_din_we),
  .iteration        (iteration),
  .first_half       (first_half),
  .first_iteration  (first_iteration),
  .cn_we            (cn_we),
  .cn_rd            (cn_rd),
  .disable_cn       (disable_cn),
  .addr_cn          (addr_cn),
  .sh_msg           (sh_msg[0]),
  .cn_msg           (cn_msg[0]),
  .dnmsg_we         (dnmsg_we_gated),
  .dnmsg_wraddr     (dnmsg_wraddr[0]),
  .dnmsg_rdaddr     (dnmsg_rdaddr[0]),
  .dnmsg_din        (dnmsg_din[0]),
  .dnmsg_dout       (dnmsg_dout[0])
);

ldpc_ram_behav #(
  .WIDTH    (17+4*(LLRWIDTH-1)+32),
  .LOG2DEPTH(7+FOLDFACTOR)
) ldpc_cnholder_0i (
  .clk(clk),
  .we(dnmsg_we_gated),
  .din(dnmsg_din[0]),
  .wraddr(dnmsg_wraddr[0]),
  .rdaddr(dnmsg_rdaddr[0]),
  .dout(dnmsg_dout[0])
);

// second - same as entire array, but is the source of the signal "we"
  ldpc_cn #( .FOLDFACTOR(FOLDFACTOR),
             .LLRWIDTH(LLRWIDTH)
  ) ldpc_cn1i(
    .clk              (clk),
    .rst              (rst),
    .llr_access       (llr_access),
    .llr_addr         (llr_addr),
    .llr_din_we       (llr_din_we),
    .iteration        (iteration),
    .first_half       (first_half),
    .first_iteration  (first_iteration),
    .cn_we            (cn_we),
    .cn_rd            (cn_rd),
    .disable_cn       (zero),
    .addr_cn          (addr_cn),
    .sh_msg           (sh_msg[1]),
    .cn_msg           (cn_msg[1]),
    .dnmsg_we         (dnmsg_we),
    .dnmsg_wraddr     (dnmsg_wraddr[1]),
    .dnmsg_rdaddr     (dnmsg_rdaddr[1]),
    .dnmsg_din        (dnmsg_din[1]),
    .dnmsg_dout       (dnmsg_dout[1])
);

  ldpc_ram_behav #(
    .WIDTH    (17+4*(LLRWIDTH-1)+32),
    .LOG2DEPTH(7+FOLDFACTOR)
  ) ldpc_cnholder_1i (
    .clk(clk),
    .we(dnmsg_we),
    .din(dnmsg_din[1]),
    .wraddr(dnmsg_wraddr[1]),
    .rdaddr(dnmsg_rdaddr[1]),
    .dout(dnmsg_dout[1])
  );

generate
  genvar k;

  for( k=2; k<NUMINSTANCES; k=k+1 )
  begin: checknodes
    ldpc_cn #( .FOLDFACTOR(FOLDFACTOR),
               .LLRWIDTH(LLRWIDTH)
    ) ldpc_cni(
      .clk              (clk),
      .rst              (rst),
      .llr_access       (llr_access),
      .llr_addr         (llr_addr),
      .llr_din_we       (llr_din_we),
      .iteration        (iteration),
      .first_half       (first_half),
      .first_iteration  (first_iteration),
      .cn_we            (cn_we),
      .cn_rd            (cn_rd),
      .disable_cn       (zero),
      .addr_cn          (addr_cn),
      .sh_msg           (sh_msg[k]),
      .cn_msg           (cn_msg[k]),
      .dnmsg_we         (),
      .dnmsg_wraddr     (dnmsg_wraddr[k]),
      .dnmsg_rdaddr     (dnmsg_rdaddr[k]),
      .dnmsg_din        (dnmsg_din[k]),
      .dnmsg_dout       (dnmsg_dout[k])
  );

    ldpc_ram_behav #(
      .WIDTH    (17+4*(LLRWIDTH-1)+32),
      .LOG2DEPTH(7+FOLDFACTOR)
    ) ldpc_cnholder_i (
      .clk(clk),
      .we(dnmsg_we),
      .din(dnmsg_din[k]),
      .wraddr(dnmsg_wraddr[k]),
      .rdaddr(dnmsg_rdaddr[k]),
      .dout(dnmsg_dout[k])
    );
  end
endgenerate

endmodule
//-------------------------------------------------------------------------
//
// File name    :  ldpc_vncluster.v
// Title        :
//              :
// Purpose      : A group of VN's and the associated RAM.  Clustering
//              : VN's around a RAM should reduce area in the ASIC
//              : implementation by using fewer, larger RAM's.  It should
//              : also ease placement by allowing placement of a number
//              : 
//
// ----------------------------------------------------------------------
// Revision History :
// ----------------------------------------------------------------------
//   Ver  :| Author   :| Mod. Date   :| Changes Made:
//   v1.0  | JTC      :| 2008/09/15  :|
// ----------------------------------------------------------------------
`timescale 1ns/10ps

module ldpc_vncluster #(
  parameter NUMVNS         = 3,
  parameter ENABLE_DISABLE = 1,
  parameter FOLDFACTOR     = 1,
  parameter LASTSHIFTWIDTH = 4,
  parameter LLRWIDTH       = 6
)(
  input clk,
  input rst,

  // LLR I/O
  input                       llr_access,
  input[7+FOLDFACTOR-1:0]     llr_addr,
  input                       llr_din_we,
  input[NUMVNS*LLRWIDTH-1:0]  llr_din,
  output[NUMVNS*LLRWIDTH-1:0] llr_dout,

  // message control
  input                   iteration,
  input                   first_half,
  input                   first_iteration,  // ignore upmsgs
  input                   we_vnmsg,
  input                   disable_vn,
  input[7+FOLDFACTOR-1:0] addr_vn,

  // message I/O
  input  wire[NUMVNS*LLRWIDTH-1:0] sh_cluster_msg,
  output wire[NUMVNS*LLRWIDTH-1:0] vn_cluster_msg
);

wire   zero;
assign zero = 0;

////////////////////////
// 2-d/1-d conversion //
////////////////////////
wire[LLRWIDTH-1:0] vn_msg[0:NUMVNS-1];
wire[LLRWIDTH-1:0] sh_msg[0:NUMVNS-1];
wire[LLRWIDTH-1:0] llr_din_2d[0:NUMVNS-1];
wire[LLRWIDTH-1:0] llr_dout_2d[0:NUMVNS-1];

generate
  genvar j;

  for( j=0; j<NUMVNS; j=j+1 )
  begin: convert1d2d
    assign vn_cluster_msg[LLRWIDTH*j+LLRWIDTH-1 -: LLRWIDTH] = vn_msg[j];
    assign sh_msg[j] = sh_cluster_msg[LLRWIDTH*j+LLRWIDTH-1 -: LLRWIDTH];
    
    assign llr_din_2d[j] = llr_din[LLRWIDTH*j+LLRWIDTH-1 -: LLRWIDTH];
    assign llr_dout[LLRWIDTH*j+LLRWIDTH-1 -: LLRWIDTH] = llr_dout_2d[j];
  end
endgenerate

//////////
// VN's //
//////////
wire                   llrram_we;
wire[7+FOLDFACTOR-1:0] vnram_wraddr;
wire[7+FOLDFACTOR-1:0] vnram_rdaddr;
wire[LLRWIDTH-1:0]     llrram_din[0:NUMVNS-1];
wire[LLRWIDTH-1:0]     llrram_dout[0:NUMVNS-1];

wire                 upmsg_we;
wire[2*LLRWIDTH+4:0] upmsg_din[0:NUMVNS-1];
wire[2*LLRWIDTH+4:0] upmsg_dout[0:NUMVNS-1];

wire upmsg_we_last;

generate
  genvar i;

  for( i=0; i<NUMVNS; i=i+1 )
  begin: varnodes
    // first
    if( i==0 )
    begin
      ldpc_vn #( .FOLDFACTOR(FOLDFACTOR),
                 .LLRWIDTH  (LLRWIDTH)
      ) ldpc_vn0i (
        .clk              (clk),
        .rst              (rst),
        .llr_access       (llr_access),
        .llr_addr         (llr_addr),
        .llr_din_we       (llr_din_we),
        .llr_din          (llr_din_2d[i]),
        .llr_dout         (llr_dout_2d[i]),
        .iteration        (iteration),
        .first_half       (first_half),
        .first_iteration  (first_iteration),
        .we_vnmsg         (we_vnmsg),
        .disable_vn(zero),
        .addr_vn          (addr_vn),
        .sh_msg           (sh_msg[i]),
        .vn_msg           (vn_msg[i]),
        .vnram_wraddr     (vnram_wraddr),
        .vnram_rdaddr     (vnram_rdaddr),
        .upmsg_we         (upmsg_we),
        .upmsg_din        (upmsg_din[i]),
        .upmsg_dout       (upmsg_dout[i])
      );
    end

    // last
    if( i==NUMVNS-1 )
    begin
      ldpc_vn #( .FOLDFACTOR(FOLDFACTOR),
                 .LLRWIDTH  (LLRWIDTH)
      ) ldpc_vnlasti (
        .clk              (clk),
        .rst              (rst),
        .llr_access       (llr_access),
        .llr_addr         (llr_addr),
        .llr_din_we       (llr_din_we),
        .llr_din          (llr_din_2d[i]),
        .llr_dout         (llr_dout_2d[i]),
        .iteration        (iteration),
        .first_half       (first_half),
        .first_iteration  (first_iteration),
        .we_vnmsg         (we_vnmsg),
        .disable_vn(disable_vn),
        .addr_vn          (addr_vn),
        .sh_msg           (sh_msg[i]),
        .vn_msg           (vn_msg[i]),
        .vnram_wraddr     (),
        .vnram_rdaddr     (),
        .upmsg_we         (upmsg_we_last),
        .upmsg_din        (upmsg_din[i]),
        .upmsg_dout       (upmsg_dout[i])
      );
    end

    if( (i!=0) && (i!=NUMVNS-1) )
    begin
      ldpc_vn #( .FOLDFACTOR(FOLDFACTOR),
                 .LLRWIDTH  (LLRWIDTH)
      ) ldpc_vni (
        .clk              (clk),
        .rst              (rst),
        .llr_access       (llr_access),
        .llr_addr         (llr_addr),
        .llr_din_we       (llr_din_we),
        .llr_din          (llr_din_2d[i]),
        .llr_dout         (llr_dout_2d[i]),
        .iteration        (iteration),
        .first_half       (first_half),
        .first_iteration  (first_iteration),
        .we_vnmsg         (we_vnmsg),
        .disable_vn(zero),
        .addr_vn          (addr_vn),
        .sh_msg           (sh_msg[i]),
        .vn_msg           (vn_msg[i]),
        .vnram_wraddr     (),
        .vnram_rdaddr     (),
        .upmsg_we         (),
        .upmsg_din        (upmsg_din[i]),
        .upmsg_dout       (upmsg_dout[i])
      );
    end
  end
endgenerate

// Combine RAM I/O's
wire[NUMVNS*(2*LLRWIDTH+5)-1:0] combined_din;
wire[NUMVNS*(2*LLRWIDTH+5)-1:0] combined_dout;

generate
  genvar k;

  for( k=0; k<NUMVNS; k=k+1 )
  begin: combine_all
    assign combined_din[k*(2*LLRWIDTH+5)+2*LLRWIDTH+4 -: 2*LLRWIDTH+5] = upmsg_din[k];
    assign upmsg_dout[k] = combined_dout[k*(2*LLRWIDTH+5)+2*LLRWIDTH+4 -: 2*LLRWIDTH+5];
  end
endgenerate

generate
  if( ENABLE_DISABLE )
  begin: split_rams
    ldpc_ram_behav #(
      .WIDTH    ((NUMVNS-1)*(2*LLRWIDTH+5)),
      .LOG2DEPTH(7+FOLDFACTOR)
    ) ldpc_vn_ram0i (
      .clk(clk),
      .we(upmsg_we),
      .din(combined_din[(NUMVNS-1)*(2*LLRWIDTH+5)-1 : 0]),
      .wraddr(vnram_wraddr),
      .rdaddr(vnram_rdaddr),
      .dout(combined_dout[(NUMVNS-1)*(2*LLRWIDTH+5)-1 : 0])
    );

    ldpc_ram_behav #(
      .WIDTH    (2*LLRWIDTH+5),
      .LOG2DEPTH(7+FOLDFACTOR)
    ) ldpc_vn_ramlasti (
      .clk(clk),
      .we(upmsg_we_last),
      .din(combined_din[NUMVNS*(2*LLRWIDTH+5)-1 -: 2*LLRWIDTH+5]),
      .wraddr(vnram_wraddr),
      .rdaddr(vnram_rdaddr),
      .dout(combined_dout[NUMVNS*(2*LLRWIDTH+5)-1 -: 2*LLRWIDTH+5])
    );
  end
  else
  begin: united_ram
    ldpc_ram_behav #(
      .WIDTH    (NUMVNS*(2*LLRWIDTH+5)),
      .LOG2DEPTH(7+FOLDFACTOR)
    ) ldpc_vn_rami (
      .clk   (clk),
      .we    (upmsg_we),
      .din   (combined_din),
      .wraddr(vnram_wraddr),
      .rdaddr(vnram_rdaddr),
      .dout  (combined_dout)
    );
  end
endgenerate

endmodule

//-------------------------------------------------------------------------
//
// File name    :  ldpc_vn.v
// Title        :
//              :
// Purpose      : Variable node holder/message calculator.  Loads llr
//              : data serially, and controls RAM's.  This module is
//              : written to be as compact as possible, since it is
//              : instantiated a large number of times.  Some outputs,
//              : especially RAM controls, are not registered.
//
// ----------------------------------------------------------------------
// Revision History :
// ----------------------------------------------------------------------
//   Ver  :| Author   :| Mod. Date   :| Changes Made:
//   v1.0  | JTC      :| 2008/07/02  :|
// ----------------------------------------------------------------------
`timescale 1ns/10ps

module ldpc_vn #(
  parameter FOLDFACTOR     = 1,
  parameter LLRWIDTH       = 6
)(
  input clk,
  input rst,

  // LLR I/O
  input                   llr_access,
  input[7+FOLDFACTOR-1:0] llr_addr,
  input                   llr_din_we,
  input[LLRWIDTH-1:0]     llr_din,
  output[LLRWIDTH-1:0]    llr_dout,

  // message control
  input                   iteration,
  input                   first_half,
  input                   first_iteration,  // ignore upmsgs
  input                   we_vnmsg,
  input                   disable_vn,
  input[7+FOLDFACTOR-1:0] addr_vn,

  // message I/O
  input[LLRWIDTH-1:0]  sh_msg,
  output[LLRWIDTH-1:0] vn_msg,

  // Attached RAM, holds iteration number, original LLR and message sum
  output[7+FOLDFACTOR-1:0] vnram_wraddr,
  output[7+FOLDFACTOR-1:0] vnram_rdaddr,
  output                   upmsg_we,
  output[2*LLRWIDTH+4:0]   upmsg_din,
  input[2*LLRWIDTH+4:0]    upmsg_dout
);

// Split RAM outputs
wire[LLRWIDTH-1:0] llr_orig;
wire[LLRWIDTH+3:0] stored_msg_sum;
wire               stored_iteration;

assign llr_orig         = upmsg_dout[LLRWIDTH-1:0];
assign stored_msg_sum   = upmsg_dout[2*LLRWIDTH+3:LLRWIDTH];
assign stored_iteration = upmsg_dout[2*LLRWIDTH+4];

/************************************************************
 * Add 1's complement numbers, assume overflow not possible *
 ************************************************************/
function[LLRWIDTH+3:0] AddNewMsg( input[LLRWIDTH+3:0] a,
                                  input[LLRWIDTH-1:0] b );
  reg               signa;
  reg               signb;
  reg[LLRWIDTH+2:0] maga;
  reg[LLRWIDTH+2:0] magb;
  
  reg[LLRWIDTH+2:0] sum;
  reg[LLRWIDTH+2:0] diffa;
  reg[LLRWIDTH+2:0] diffb;
  
  reg               add;
  reg               b_big;
  reg               sign;
  reg[LLRWIDTH+3:0] result;
  
begin
  // strip out magnitude and sign bits
  signa = a[LLRWIDTH+3];
  signb = b[LLRWIDTH-1];
  maga  = a[LLRWIDTH+2:0];
  magb  = { 4'b0000, b[LLRWIDTH-2:0] };

  // basic calculations
  sum   = maga + magb;
  diffa = maga - magb;
  diffb = magb - maga;
  
  // control bits
  add   = signa==signb;
  b_big = maga<magb;
  sign  = b_big ? signb : signa;

  if( add )
    result = { sign, sum };
  else if( b_big )
    result = { sign, diffb };
  else
    result = { sign, diffa };

  AddNewMsg = result;
end
endfunction

/*************************************************
 * Saturate message to fewer bits before passing *
 *************************************************/
function[LLRWIDTH-1:0] SaturateMsg( input[LLRWIDTH+3:0] a );
begin
  if( a[LLRWIDTH+2:LLRWIDTH-1] != 4'b0000 )
    SaturateMsg[LLRWIDTH-2:0] = { (LLRWIDTH-1){1'b1} };
  else
    SaturateMsg[LLRWIDTH-2:0] = a[LLRWIDTH-2:0];
  
  SaturateMsg[LLRWIDTH-1] = a[LLRWIDTH+3];
end
endfunction

/********************************************
 * Delays to align controls with RAM output *
 ********************************************/
localparam RAM_LATENCY = 2;

integer loopvar1;

reg[7+FOLDFACTOR-1:0] vnram_rdaddr_int;

reg[LLRWIDTH-1:0]     sh_msg_del[0:RAM_LATENCY-1];
reg                   we_vnmsg_del[0:RAM_LATENCY-1];
reg[7+FOLDFACTOR-1:0] vnram_rdaddr_del[0:RAM_LATENCY-1];
reg                   disable_del[0:RAM_LATENCY-1];    

wire[LLRWIDTH-1:0]     sh_msg_aligned_ram;
wire                   we_vnmsg_aligned_ram;
wire[7+FOLDFACTOR-1:0] vnram_rdaddr_aligned_ram;
wire                   disable_aligned_ram;

reg recycle_result;

// mux in alternative address for final read-out
assign vnram_rdaddr = vnram_rdaddr_int;
always @( * ) vnram_rdaddr_int <= #1 llr_access ? llr_addr : addr_vn;

assign sh_msg_aligned_ram       = sh_msg_del[RAM_LATENCY-1];
assign we_vnmsg_aligned_ram     = we_vnmsg_del[RAM_LATENCY-1];
assign vnram_rdaddr_aligned_ram = vnram_rdaddr_del[RAM_LATENCY-1];
assign disable_aligned_ram      = disable_del[RAM_LATENCY-1];    

always @( posedge rst, posedge clk )
  if( rst )
  begin
    for( loopvar1=0; loopvar1<RAM_LATENCY; loopvar1=loopvar1+1 )
    begin
      sh_msg_del[loopvar1]       <= 0;
      we_vnmsg_del[loopvar1]     <= 0;
      vnram_rdaddr_del[loopvar1] <= 0;
      disable_del[loopvar1]      <= 0;
    end
    recycle_result <= 0;
  end
  else
  begin
    sh_msg_del[0]        <= sh_msg;
    we_vnmsg_del[0]      <= we_vnmsg;
    vnram_rdaddr_del[0]  <= vnram_rdaddr_int; 
    disable_del[0]       <= disable_vn;

    for( loopvar1=1; loopvar1<RAM_LATENCY; loopvar1=loopvar1+1 )
    begin
      sh_msg_del[loopvar1]       <= sh_msg_del[loopvar1 -1];
      we_vnmsg_del[loopvar1]     <= we_vnmsg_del[loopvar1 -1];
      vnram_rdaddr_del[loopvar1] <= vnram_rdaddr_del[loopvar1 -1];
      disable_del[loopvar1]      <= disable_del[loopvar1 -1];
    end
    
    // Use previous result rather than the RAM contents for two adjacent
    // writes to the same address
    recycle_result <= (vnram_rdaddr_aligned_ram==vnram_rdaddr_del[RAM_LATENCY-2]) &
                      we_vnmsg_aligned_ram & we_vnmsg_del[RAM_LATENCY-2];
  end

/************************
 * Message calculations *
 ************************/
// Add initial LLR to message offset (except for first iteration)
reg[LLRWIDTH+3:0]  msg0_norst;
wire[LLRWIDTH+3:0] msg0;
reg[LLRWIDTH-1:0]  msg1;

wire start_new_upmsg;
reg  rst_msg0;

wire[LLRWIDTH+3:0] msg_sum;

reg[LLRWIDTH+3:0] msg_sum_reg;

// Add upmsg to the result, except:
// - during first iteration, since no upmsg exists
// - first message of each new iteration, where upmsg needs to be reset
assign start_new_upmsg = (stored_iteration!=iteration) & we_vnmsg_aligned_ram;

assign msg0 = rst_msg0 ? 0 : msg0_norst;

always @( posedge clk, posedge rst )
  if( rst )
  begin
    msg0_norst  <= 0;
    rst_msg0    <= 0;
    msg1        <= 0;
    msg_sum_reg <= 0;
  end
  else
  begin
    // msg0 = sum of received upstream messages
    // clear msg0 when beginning a new set of upstream messages
    msg0_norst <= recycle_result ? msg_sum : stored_msg_sum;
    rst_msg0   <= start_new_upmsg & ~recycle_result;
    
    msg1 <= (llr_access || first_half) ? llr_orig : sh_msg_aligned_ram;
    
    msg_sum_reg <= msg_sum;
  end

// When creating downstream messages, or preparing final result:
//      msg_sum = llr + sum of messages
// When receiving upstream messages:
//      msg_sum = new message + sum of messages
assign msg_sum = AddNewMsg( msg0, msg1 );

/****************************************
 * Delay controls to align with msg_sum *
 ****************************************/
localparam CALC_LATENCY = 2;

integer loopvar2;

reg                   we_vnmsg_del2[0:RAM_LATENCY-1];
reg[7+FOLDFACTOR-1:0] vnram_rdaddr_del2[0:RAM_LATENCY-1];
reg[LLRWIDTH-1:0]     llrram_dout_del2[0:RAM_LATENCY-1];
reg                   disable_del2[0:RAM_LATENCY-1];    

wire                   we_vnmsg_aligned_msg;
wire[7+FOLDFACTOR-1:0] vnram_rdaddr_aligned_msg;
wire[LLRWIDTH-1:0]     llrram_dout_aligned_msg;
wire                   disable_aligned_msg;

assign we_vnmsg_aligned_msg     = we_vnmsg_del2[RAM_LATENCY-1];
assign vnram_rdaddr_aligned_msg = vnram_rdaddr_del2[RAM_LATENCY-1];
assign llrram_dout_aligned_msg  = llrram_dout_del2[RAM_LATENCY-1];
assign disable_aligned_msg      = disable_del2[RAM_LATENCY-1];    

always @( posedge rst, posedge clk )
  if( rst )
  begin
    for( loopvar2=0; loopvar2<RAM_LATENCY; loopvar2=loopvar2+1 )
    begin
      we_vnmsg_del2[loopvar2]     <= 0;
      vnram_rdaddr_del2[loopvar2] <= 0;
      llrram_dout_del2[loopvar2]  <= 0;
      disable_del2[loopvar2]      <= 0;
    end
  end
  else
  begin
    we_vnmsg_del2[0]      <= we_vnmsg_aligned_ram;
    vnram_rdaddr_del2[0]  <= vnram_rdaddr_aligned_ram; 
    llrram_dout_del2[0]   <= llr_orig;
    disable_del2[0]       <= disable_aligned_ram;

    for( loopvar2=1; loopvar2<RAM_LATENCY; loopvar2=loopvar2+1 )
    begin
      we_vnmsg_del2[loopvar2]     <= we_vnmsg_del2[loopvar2 -1];
      vnram_rdaddr_del2[loopvar2] <= vnram_rdaddr_del2[loopvar2 -1];
      llrram_dout_del2[loopvar2]  <= llrram_dout_del2[loopvar2 -1];
      disable_del2[loopvar2]      <= disable_del2[loopvar2 -1];
    end
  end

/*******************************
 * Write message totals to RAM *
 *******************************/
reg[7+FOLDFACTOR-1:0] vnram_wraddr_int;
reg[LLRWIDTH-1:0]     new_llr;
reg                   new_iteration;
reg[LLRWIDTH+3:0]     new_msg_sum;
reg                   upmsg_we_int;

assign vnram_wraddr = vnram_wraddr_int;
assign upmsg_din    = { new_iteration, new_msg_sum, new_llr };
assign upmsg_we     = upmsg_we_int;

always @( posedge rst, posedge clk )
  if( rst )
  begin
    vnram_wraddr_int <= 0;
    new_llr          <= 0;
    new_msg_sum      <= 0;
    new_iteration    <= 0;
    upmsg_we_int     <= 1;
  end
  else
  begin
    // mux and register outputs
    vnram_wraddr_int <= #1 llr_access ? llr_addr : vnram_rdaddr_aligned_msg;
    new_llr          <= #1 llr_access ? llr_din  : llrram_dout_aligned_msg;
    new_msg_sum      <= #1 llr_access ? 0        : msg_sum_reg;
    
    new_iteration    <= #1 llr_access | iteration;
    
    upmsg_we_int     <= #1 ~(llr_din_we | (we_vnmsg_aligned_msg & ~disable_aligned_msg));
  end

/*****************************************************************
 * Saturate message to fewer bits for message passing and output *
 *****************************************************************/
reg[LLRWIDTH-1:0] vn_msg_int;

assign llr_dout = vn_msg_int;
assign vn_msg   = vn_msg_int;

always @( posedge rst, posedge clk )
  if( rst )
    vn_msg_int <= 0;
  else
    vn_msg_int <= SaturateMsg(msg_sum_reg);

endmodule

